!VERSION:  17_03
!AUTHORS:  C1-C3   Burcat   
!NOTE:     SPECIES RE-ARRANGED AS THE SAME ORDER IN MECH
!
!VERSION:  17_05
!Following species are updated from Burcat's Database:Kik
! C6H5CHCH3	FLUORENE	C5H6	INDENYL	C14H19	C12H7	C12H9        
! C6H5CH2C6H5	C10H7	CH3C6H4	C6H5C2H	C6H5O	C6H5C2H3	C10H7CH3
! C10H7CHO	RXYLENE	C10H7CH2	XYLENE	C6H2	Toluene	C6H5OH
! C14H10	C6H5C2H4C6H5	C4H2	C16H10	C5H5CH3	C7H7	BENZYNE
! C6H5C2H2	C12H8	C6H5C2H5	C10H7O	BENZENE	C4H4	INDENE
! C5H5	C10H6CH3	C6H5 	C10H8	FULVENE	BIPHENYL	C6H4C2H
!Following species are updated from ATcT's Database:Ghobad
! H	H2	O	O2	HE
! OH	H2O	N2	HO2	HCO
! H2O2	AR	CO	CO2

THERMO
300.   1000.   4000.
!Work C5
cC7H7 Cyheptatrie A09/05C  7.H  7.   0.   0.G   200.000  6000.000 1000.        1
 1.37839351E+01 2.32922891E-02-8.36543230E-06 1.35064040E-09-8.08726926E-14    2
 2.71779724E+04-4.85624908E+01 1.37723080E+00 3.27432725E-02 4.58225372E-05    3
-9.07721756E-08 4.08096948E-11 3.16491191E+04 2.10799820E+01 3.37597997E+04    4
A1C7              T 7/98C  11H   9    0    0G   200.000  6000.000 1000.        1 ! methyl naphthalene Burcat kik 1-C10H7-CH2*
 2.18977539E+01 3.26102636E-02-1.18401218E-05 1.92574628E-09-1.15903442E-13    2
 2.24571098E+04-9.41050741E+01-2.53234304E+00 7.32920338E-02 2.02974707E-05    3
-9.36547823E-08 4.70753594E-11 3.02906705E+04 3.79638513E+01 3.28097266E+04    4
! From Marco  RF
DECA_ET                 C  10H  16O   1    0G   300.000  5000.000 1425.000    01
 2.93462856E+01 4.07923202E-02-1.37934492E-05 2.12631155E-09-1.22794883E-13    2
-4.03406303E+04-1.40206695E+02-2.78036486E+01 1.90456576E-01-1.63231397E-04    3
 6.93353094E-08-1.15568584E-11-2.25640096E+04 1.60227296E+02                   4
C10H16                  C  10H  16    0    0G   300.000  5000.000 1383.000    01
 3.00622157E+01 4.04814732E-02-1.43100916E-05 2.27150755E-09-1.33848364E-13    2
-2.64487109E+04-1.50795570E+02-1.59752190E+01 1.41881956E-01-9.68191663E-05    3
 3.15855617E-08-3.94115263E-12-9.95822808E+03 9.84523499E+01                   4
C10H15                  C  10H  15    0    0G   300.000  5000.000 1388.000    01
 3.06775047E+01 3.73366921E-02-1.32088842E-05 2.09790798E-09-1.23671129E-13    2
-8.63138773E+03-1.55587564E+02-1.68540337E+01 1.46145526E-01-1.06465345E-04    3
 3.76155230E-08-5.19112395E-12 7.91843171E+03 1.00180731E+02                   4
C6H5C4H9      3/99      C  10H  14    0    0G   300.000  5000.000 1395.000    41
 2.67352334E+01 3.43477266E-02-1.17087252E-05 1.81434544E-09-1.05143951E-13    2
-1.51216286E+04-1.18171023E+02-6.22856223E+00 1.13691752E-01-8.50361112E-05    3
 3.27496505E-08-5.12339478E-12-3.97172741E+03 5.79294597E+01                   4
RC6H5C4H8     3/99      C  10H  130   00   0G   300.000  5000.000 1393.000    41
 2.70273993E+01 3.21704122E-02-1.10893400E-05 1.73097280E-09-1.00815459E-13    2
 2.35147019E+03-1.20696474E+02-3.97290080E+00 1.05990334E-01-7.87536684E-05    3
 3.01569625E-08-4.71350779E-12 1.29600077E+04 4.52696443E+01                   4
C6H5C4H7-3    8/99 THERMC  10H  12    0    0G   300.000  5000.000 1395.000    31  !TETRALIN
 2.53129170E+01 3.14281387E-02-1.08152689E-05 1.68620292E-09-9.81246226E-14    2
-1.40337072E+03-1.10601858E+02-5.52864894E+00 1.07276062E-01-8.33212344E-05    3
 3.36538598E-08-5.55115817E-12 8.92646491E+03 5.36875671E+01                   4
RC6H5C4H8OO  21/13 THERMC  10H  13O   2    0G   300.000  5000.000 1384.000    61
 3.29433924E+01 3.24682623E-02-1.24870478E-05 2.07708155E-09-1.25876772E-13    2
-1.26391156E+04-1.46881012E+02-3.28758026E+00 1.13009541E-01-8.07422394E-05    3
 2.85337544E-08-4.11461923E-12 4.66204317E+02 4.93485667E+01                   4
QC6H5C4H8     6/ 3/99   C  10H  13O   2    0G   300.000  5000.000 1391.000    61
 3.18818252E+01 3.27029227E-02-1.13668697E-05 1.78433731E-09-1.04337691E-13    2
-5.51050095E+03-1.36501133E+02-4.64927400E+00 1.21423535E-01-9.46502187E-05    3
 3.77087559E-08-6.09386626E-12 6.80419866E+03 5.84407930E+01                   4
QC6H5C4H8OO        THERMC  10H  13O   4    0G   300.000  5000.000 1394.000    71
 3.61027915E+01 3.40077547E-02-1.18624314E-05 1.86619563E-09-1.09279047E-13    2
-2.54960378E+04-1.55903949E+02-3.49701990E+00 1.36010314E-01-1.15199287E-04    3
 5.03824666E-08-8.90327014E-12-1.26357910E+04 5.35021839E+01                   4
KETBBZ         99 THERM C  10H  12O   3    0G   300.000  5000.000 1391.000    61
 3.36726156E+01 3.15259909E-02-1.10345070E-05 1.73992324E-09-1.02047241E-13    2
-1.33627844E+04-1.46053045E+02-2.68620243E+00 1.23388659E-01-1.02246011E-04    3
 4.37989670E-08-7.61792966E-12-1.36674405E+03 4.68663270E+01                   4
IC12-OQOOH              C  12H  24O   3     G    300.00   4000.00 1678.00      1
 .447068212E+02 .522272795E-01-.195350799E-04 .322923457E-08-.195935332E-12    2
-.818914807E+05-.192299360E+03 .877388676E+01 .119113497E+00-.561329021E-04    3
 .677643630E-08 .106366869E-11-.685051188E+05 .572134782E+01                   4
IC12H26                 C  12H  26          G    300.00   4000.00 1391.00      1
 .385099212E+02 .563550048E-01-.191493200E-04 .296024862E-08-.171244150E-12    2
-.548849270E+05-.169785166E+03-.262181594E+01 .147237711E+00-.943970271E-04    3
 .307441268E-07-.403602230E-11-.400654253E+05 .529882396E+02                   4
RODECOO                 C  10H  17O   2     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
QODECOOH                C  10H  17O   2     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
IC12H25                 C  12H  25          G    300.00   4000.00 1387.00      1
 .379559371E+02 .541231481E-01-.184408520E-04 .285618139E-08-.165452331E-12    2
-.312698454E+05-.166157365E+03-.117025753E+01 .136564242E+00-.813840519E-04    3
 .231564976E-07-.240764498E-11-.167979250E+05 .471339366E+02                   4
IC12-QOOH               C  12H  25O   2     G    300.00   4000.00 1392.00      1
 .427882927E+02 .547351985E-01-.185693137E-04 .286771608E-08-.165782124E-12    2
-.451897912E+05-.183774591E+03 .457142729E+00 .149660990E+00-.984019129E-04    3
 .327982507E-07-.438634589E-11-.301386488E+05 .448987214E+02                   4
IC12H25-OO              C  12H  25O   2     G    300.00   4000.00 1392.00      1
 .410672882E+02 .571682582E-01-.196096581E-04 .304996352E-08-.177163659E-12    2
-.498119415E+05-.176403781E+03 .761653139E+00 .147870053E+00-.980093227E-04    3
 .342486611E-07-.502171364E-11-.353144020E+05 .415448990E+02                   4
IC12-OOQOOH             C  12H  25O   4     G    300.00   4000.00 1393.00      1
 .478223133E+02 .563342752E-01-.193784199E-04 .302016363E-08-.175696376E-12    2
-.648031378E+05-.208209874E+03 .250560092E+01 .157994999E+00-.105503812E-03    3
 .358709948E-07-.494871123E-11-.486270464E+05 .366890378E+02                   4
! End of From Marco
! From PAH 1906 
C6H5C2H4 A1CH2CH2* 11/04C  8.H  9.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik. ER add this species in PAH1906
 1.61326962E+01 2.82904273E-02-1.01801876E-05 1.64176637E-09-9.81375329E-14    2
 2.08791061E+04-6.00115413E+01 7.33299107E-01 4.59053158E-02 3.78257231E-05    3
-9.12367411E-08 4.25589678E-11 2.61572945E+04 2.50411074E+01 2.85902549E+04    4
C18H14 C9H7C9H7         H  14C  18          G   100.000  5000.000  990.27      1  !Kik add from Jin Hanfeng Combustion and Flame 206 (2019): 1-20.
 3.20125595E+01 5.89532847E-02-2.32102353E-05 4.57752278E-09-3.44228657E-13    2
 2.23209936E+04-1.51408560E+02-1.99662811E+00 8.71499057E-02 9.94525782E-05    3
-1.89332690E-07 7.67158406E-11 3.44098058E+04 3.93622783E+01                   4
! End of  PAH 1906 

CH2OHCOOH               C   2H   4O   3     G    200.00   6000.00 1000.00      1   ! Burcat
 1.27662941E+01 1.02143437E-02-3.63547001E-06 5.83491588E-10-3.47179974E-14    2
-7.53528536E+04-3.96511752E+01 2.80443702E+00 2.10851644E-02 3.35863233E-05    3
-7.02669107E-08 3.26849274E-11-7.20649998E+04 1.51180675E+01-7.01183834E+04    4
CHOHCO2H2              C   2H   3O   3     G    200.00   6000.00 1000.00       1    !Burcat  - taken from another isomer; if = reactions present: TO BE REVISED
 1.27662941E+01 1.02143437E-02-3.63547001E-06 5.83491588E-10-3.47179974E-14    2
-7.53528536E+04-3.96511752E+01 2.80443702E+00 2.10851644E-02 3.35863233E-05    3
-7.02669107E-08 3.26849274E-11-7.20649998E+04 1.51180675E+01-7.01183834E+04    4
CHOHCO                 C   2H   4O   3     G    200.00   6000.00 1000.00       1   ! Burcat
 7.25265886E+00 7.09713194E-03-2.49703662E-06 3.97702132E-10-2.35907799E-14    2
-2.14840657E+04-9.51330315E+00 3.35107651E+00 1.55375306E-02-4.45397177E-06    3
-6.25820983E-09 4.05044001E-12-2.03011991E+04 1.11760714E+01-1.86612868E+04    4
CH3CH2COOH             C   3H   6O   2     G    200.00   6000.00 1000.00       1    !Burcat
 1.27662941E+01 1.02143437E-02-3.63547001E-06 5.83491588E-10-3.47179974E-14    2
-7.53528536E+04-3.96511752E+01 2.80443702E+00 2.10851644E-02 3.35863233E-05    3
-7.02669107E-08 3.26849274E-11-7.20649998E+04 1.51180675E+01-7.01183834E+04    4 
CH3CHCO2H2             C   3H   6O   2     G    200.00   6000.00 1000.00       1    !Burcat - taken from another isomer; if = reactions present: TO BE REVISED
 1.27662941E+01 1.02143437E-02-3.63547001E-06 5.83491588E-10-3.47179974E-14    2
-7.53528536E+04-3.96511752E+01 2.80443702E+00 2.10851644E-02 3.35863233E-05    3
-7.02669107E-08 3.26849274E-11-7.20649998E+04 1.51180675E+01-7.01183834E+04    4 
QPENTANOIC              C   5H   9O   4     G    300.00   4000.00 1386.00      1    !taken from alcohol they don't matter as Lumped
 .129455763E+02 .795235476E-02-.280679691E-05 .445205248E-09-.262240810E-13    2
 .175946397E+05-.478819894E+02-.584674088E+01 .620875882E-01-.630010605E-04    3
 .306882361E-07-.575456234E-11 .230253176E+05 .492940922E+02                   4
RO2PENTANOIC            C   5H   9O   4     G    300.00   4000.00 1392.00      1     !taken from alcohol they don't matter as Lumped
 .179101133E+02 .211247449E-01-.724787505E-05 .112742547E-08-.654930094E-13    2
-.371878276E+05-.612769774E+02 .289779336E+01 .560720331E-01-.390996379E-04    3
 .147174953E-07-.234862827E-11-.318812119E+05 .195265598E+02                   4
ZPENTANOIC              C   5H   9O   6     G    300.00   4000.00 1397.00      1      !taken from alcohol they don't matter as Lumped
 .236719411E+02 .205751255E-01-.708127339E-05 .110392970E-08-.642301320E-13    2
-.515463449E+05-.860806755E+02 .475209184E+01 .678608013E-01-.534336966E-04    3
 .221852722E-07-.378003417E-11-.452511232E+05 .144907043E+02                   4
KPENTANOIC              C   5H   8O   5     G    300.00   4000.00 1396.00      1        !taken from alcohol they don't matter as Lumped
 .219367270E+02 .180406285E-01-.626171080E-05 .981855896E-09-.573639516E-13    2
-.664546784E+05-.813588272E+02-.445736457E+01 .947202096E-01-.937478682E-04    3
 .464802131E-07-.899314409E-11-.587131282E+05 .551970961E+02                   4
QBUTANOIC               C   4H   7O   4     G    300.00   4000.00 1386.00      1    !taken from alcohol they don't matter as Lumped
 .129455763E+02 .795235476E-02-.280679691E-05 .445205248E-09-.262240810E-13    2
 .175946397E+05-.478819894E+02-.584674088E+01 .620875882E-01-.630010605E-04    3
 .306882361E-07-.575456234E-11 .230253176E+05 .492940922E+02                   4
RO2BUTANOIC             C   4H   7O   4     G    300.00   4000.00 1392.00      1     !taken from alcohol they don't matter as Lumped
 .179101133E+02 .211247449E-01-.724787505E-05 .112742547E-08-.654930094E-13    2
-.371878276E+05-.612769774E+02 .289779336E+01 .560720331E-01-.390996379E-04    3
 .147174953E-07-.234862827E-11-.318812119E+05 .195265598E+02                   4
ZBUTANOIC               C   4H   7O   6     G    300.00   4000.00 1397.00      1      !taken from alcohol they don't matter as Lumped
 .236719411E+02 .205751255E-01-.708127339E-05 .110392970E-08-.642301320E-13    2
-.515463449E+05-.860806755E+02 .475209184E+01 .678608013E-01-.534336966E-04    3
 .221852722E-07-.378003417E-11-.452511232E+05 .144907043E+02                   4
KBUTANOIC               C   4H   6O   5     G    300.00   4000.00 1396.00      1        !taken from alcohol they don't matter as Lumped
 .219367270E+02 .180406285E-01-.626171080E-05 .981855896E-09-.573639516E-13    2
-.664546784E+05-.813588272E+02-.445736457E+01 .947202096E-01-.937478682E-04    3
 .464802131E-07-.899314409E-11-.587131282E+05 .551970961E+02                   4
CYC5H4CO                C   6H   4O   1     G    300.00   4000.00 1000.00      1   ! molecola da furutani 2017 calcolare termo con automech
 .137221720E+02 .174688771E-01-.635504520E-05 .103492308E-08-.623410504E-13    2
 15.2872748E+03-.488181680E+02-.466204455E+00 .413443975E-01 .132412991E-04    3
-.572872769E-07 .289763707E-10 1.97785839E+04 .276990274E+02                   4
C6H4O                   C   6H   4O   1     G    300.00   4000.00 1000.00      1   ! Biradicale da guaiacolo rivedeer sono quelle di C6H5O
 .137221720E+02 .174688771E-01-.635504520E-05 .103492308E-08-.623410504E-13    2
 15.2872748E+03-.488181680E+02-.466204455E+00 .413443975E-01 .132412991E-04    3
-.572872769E-07 .289763707E-10 1.97785839E+04 .276990274E+02                   4
!RPHENPH                 C   6H   5O   1     G    300      3500    1000         1
! 7.48628748E+00 3.11726354E-02-1.63674822E-05 4.10796074E-09-3.98797024E-13    2    
! 1.49961514E+04-1.26543728E+01-8.11677970E+00 9.35849042E-02-1.09985886E-04    3    
! 6.65202295E-08-1.60018642E-11 1.81167649E+04 6.26214070E+01                   4    
RCATEPH                 C   6H   5O   2     G    300      3500    1000         1
 1.18218904E+01 2.70911132E-02-1.34162451E-05 3.08575091E-09-2.72411991E-13    2    
-7.82412443E+03-3.10506043E+01-7.41421113E+00 1.04035520E-01-1.28832855E-04    3    
 8.00301573E-08-1.95085136E-11-3.97690414E+03 6.17524664E+01                   4    
C6H4C2H3          T12/07C  8.H  7.   0.   0.G   200.000  6000.000 1000.00      1
 1.57334515E+01 2.38965492E-02-8.60829763E-06 1.39223384E-09-8.35065775E-14    2
 4.08827573E+04-5.82476667E+01 1.17830774E+00 3.40765502E-02 5.85065530E-05    3
-1.10953244E-07 4.95222636E-11 4.61414992E+04 2.36053284E+01 4.83284254E+04    4
C7H6O3                  C   7H   6O   3     G    300      3500    1000         1
 9.6100307E+00  4.6312670E-02 -2.4985466E-05  6.2313178E-09 -5.9678291E-13     2
-5.2881308E+04 -1.4662558E+01 -7.0701097E+00  1.1303323E-01 -1.2506631E-04     3
 7.2951879E-08 -1.7276923E-11 -4.9545280E+04  6.5809478E+01                    4
RC7H5O3                 C   7H   5O   3     G    300      3500    1000         1
 1.03519980E+01 4.06949717E-02-2.16398081E-05 5.16863129E-09-4.69580170E-13    2
-3.48541024E+04-1.78724727E+01-6.94106227E+00 1.09867214E-01-1.25398170E-04    3
 7.43408724E-08-1.77626405E-11-3.13954904E+04 6.55565469E+01                   4
C8H6O3                  C   8H   6O   3     G    300      3500    1000         1
 4.593105E+00   6.232992E-02  -3.473750E-05   8.749391E-09  -8.397915E-13      2
-4.481918E+04   1.511354E+01  -8.470549E+00   1.145845E-01  -1.131194E-04      3
 6.100401E-08  -1.390345E-11  -4.220645E+04   7.813812E+01                     4
RGUAIPH                 C   7H   7O   2     G    300      3500    1000         1
 1.0328870E+01  4.1581495E-02 -2.2022073E-05  5.3914934E-09 -5.0157294E-13     2
-4.9145545E+03 -2.2004822E+01 -7.2388396E+00  1.1185234E-01 -1.2742833E-04     3
 7.5662334E-08 -1.8069283E-11 -1.4010125E+03  6.2749224E+01                    4
RSALICPH                C   7H   5O   2     G    300      3500    1000         1
 6.006532E+00   4.553370E-02  -2.518536E-05   6.391630E-09  -6.195741E-13      2
 4.679999E+02   2.823677E+00  -8.006329E+00   1.015851E-01  -1.092625E-04      3
 6.244307E-08  -1.463244E-11   3.270572E+03   7.042763E+01                     4
C6H4OCH3                C   7H   7O   1     G    300      3500    1000         1
 6.1403860E+00  4.5274166E-02 -2.4649522E-05  6.3063297E-09 -6.1560301E-13     2
 1.7881392E+04 -4.3538799E+00 -8.0284207E+00  1.0194939E-01 -1.0966236E-04     3
 6.2981557E-08 -1.4784410E-11  2.0715154E+04  6.4002422E+01                    4
CATECHOL                C   6H   6O   2     G    300.00   3500.00 1150.00      1
 1.43499796e+01 2.44086040e-02-1.04210961e-05 2.01938934e-09-1.47232776e-13    2
-3.94515398e+04-4.76262851e+01-5.49815264e+00 9.34455856e-02-1.00469333e-04    3
 5.42212658e-08-1.14954668e-11-3.48864694e+04 5.09034930e+01                   4
OC6H4OH                 C   6H   5O   2     G    300.00   3500.00 1140.00      1
 1.40810368e+01 2.16036559e-02-9.34848731e-06 1.81734390e-09-1.31737736e-13    2
-2.57458617e+04-4.55416672e+01-4.82568614e+00 8.79430347e-02-9.66371436e-05    3
 5.28633417e-08-1.13260355e-11-2.14351289e+04 4.81496570e+01                   4
OC6H4OH                 H  5 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! DHof -32.74 O-OC6H4OH W13 LPM automech from C6H5+O2 paper
 9.05445252E+00 3.27089888E-02-1.69405687E-05 4.23212572E-09-4.13426536E-13    2
-2.34445619E+04-2.26110686E+01-1.57606826E-02 4.37516112E-02 1.47150643E-05    3
-5.88273942E-08 2.90180512E-11-2.05689532E+04 2.68352761E+01                   4
P-OC6H4OH               H  5 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! DHof -26.91 W16, NOT IN FINAL LUMPED MECH
 1.04799021E+01 3.06270960E-02-1.59736238E-05 4.01775452E-09-3.94850716E-13    2
-2.08131901E+04-2.97663019E+01 6.87475479E-02 4.72745543E-02 5.84712321E-06    3
-5.06271974E-08 2.61930505E-11-1.76556892E+04 2.61615828E+01                   4
O-C6H4O2H               H  5 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! DHof -11.77 LPM automech from C6H5+O2 paper
 8.68756237E+00 3.37206762E-02-1.76439955E-05 4.43399930E-09-4.34621804E-13    2
-1.25169228E+04-1.76564145E+01 1.37781528E+00 3.99178050E-02 1.67600872E-05    3
-5.63411958E-08 2.70491089E-11-1.00767150E+04 2.28258250E+01                   4
GUAIACOL                C   7H   8O   2     G    300.00   3500.00 1000.00      1
 9.99301751e+00 4.50609491e-02-2.36180835e-05 5.74985960e-09-5.33615080e-13    2
-3.55531886e+04-2.30989118e+01-7.52910597e+00 1.15149443e-01-1.28750824e-04    3
7.58383535e-08 -1.80557386e-11-3.20487639e+04 6.14352053e+01                   4
SALICALD                C   7H   6O   2     G    300.00   3500.00 1000.00      1
 1.64419508E+01 2.56565170E-02-9.29837990E-06 1.30953013E-09-5.02395383E-14    2
-3.38514104E+04-5.63974383E+01-4.36490575E-01 5.47073717E-02-7.07267500E-07    3
-3.69175398E-08 1.74133046E-11-2.82980420E+04 3.52247637E+01                   4
VANILLIN                C   8H   8O   3     G    300.00   3500.00 1260.00      1
 1.36544650e+01 4.84143232e-02-2.42641798e-05 5.50487829e-09-4.76001947e-13    2
-5.18855416e+04-3.54575728e+01-4.86637458e+00 1.07210639e-01-9.42597942e-05    3
 4.25395949e-08-7.82416000e-12-4.72182900e+04 5.81751551e+01                   4
!   ---------ARAMCO 2.0 -------------------
C3H6       8/12/15      C   3H   6    0    0G   298.000  6000.000 1000.000    01
 6.59032304E+00 1.52592866E-02-5.30369441E-06 8.35510888E-10-4.91215549E-14    2
-2.47481113E+02-1.15748238E+01-1.54606737E+00 4.36553128E-02-5.61392417E-05    3
 4.98421927E-08-1.84798923E-11 2.07056233E+03 2.99232495E+01                   4
C3H5-A     8/12/15      C   3H   5    0    0G   298.000  6000.000 1000.000    01
 7.37604097E+00 1.23449782E-02-4.26463882E-06 6.69045835E-10-3.92202554E-14    2
 1.77332960E+04-1.61758204E+01-3.32899442E+00 5.38423469E-02-7.65500752E-05    3
 6.35512285E-08-2.14283003E-11 2.03420628E+04 3.68038362E+01                   4
C3H5-S     8/12/15      C   3H   5    0    0G   300.000  5000.000 1390.000    11
 7.95954498E+00 1.11163183E-02-3.75197834E-06 5.77246260E-10-3.32768957E-14    2
 2.80567891E+04-1.79800372E+01 1.61793372E+00 2.44803904E-02-1.41856503E-05    3
 4.16402233E-09-4.90904795E-13 3.04291037E+04 1.66341443E+01                   4
C3H5-T     8/12/15      C   3H   5    0    0G   300.000  5000.000 1376.000    11
 7.69949212E+00 1.17803985E-02-4.07791749E-06 6.38119222E-10-3.72229675E-14    2
 2.61747145E+04-1.68305890E+01 2.29256998E+00 1.98527646E-02-6.42635654E-06    3
-5.90016395E-10 5.05491095E-13 2.85773377E+04 1.39407124E+01                   4
!   --------- end ARAMCO 2.0 -------------------
LC5H8                   C   5H   8          G    300.00   4000.00 1000.00      1
 .797205310E+01 .268614160E-01-.956546320E-05 .113079120E-08 .000000000E+00    2
 .510466811E+04-.185090870E+02 .176636500E+01 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .684030700E+04 .137180600E+02                   4
CYC5H8                  C   5H   8          G    300.00   4000.00 1000.00      1
 .772447728E+01 .283223160E-01-.115452360E-04 .215408150E-08-.150541780E-12    2
-.782614232E+03-.197696844E+02 .268981400E+01 .209545500E-02 .113036870E-03    3
-.154080700E-06 .627636580E-10 .231396630E+04 .152940560E+02                   4
CYC6H8                  C   6H   8          G    300.00   4000.00 1384.00      1
 .167797183E+02 .200748305E-01-.710732570E-05 .112925397E-08-.665827513E-13    2
 .222453062E+04-.729120687E+02-.719572313E+01 .780676798E-01-.620002183E-04    3
 .253310854E-07-.423684696E-11 .104082650E+05 .552451233E+02                   4
CYC6H10                 C   6H  10          G    300.00   4000.00 1388.00      1
 .164687940E+02 .250464584E-01-.873323457E-05 .137353265E-08-.804138942E-13    2
-.977694533E+04-.696690108E+02-.607599781E+01 .751138370E-01-.506516889E-04    3
 .171683701E-07-.235089637E-11-.166592755E+04 .523699408E+02                   4
DIALLYL                 C   6H  10          G    300.00   4000.00 1413.00      1
 .160456030E+02 .234774145E-01-.785797929E-05 .120200542E-08-.690100029E-13    2
 .211899382E+04-.588452460E+02-.101375402E+01 .638242808E-01-.440653860E-04    3
 .158295163E-07-.230830701E-11 .794033696E+04 .325056094E+02                   4
LC5H7 1,4diene-3ylA 1/05C  5.H  7.   0.   0.G   200.000  6000.000 1000.        1      ! CVCCJCVC in itvcreck, but wrong thermodynamics
 1.01206141E+01 2.19623708E-02-8.13808356E-06 1.32677709E-09-7.97014062E-14    2
 1.97304588E+04-2.73862410E+01 2.36470149E+00 2.39388874E-02 3.85164588E-05    3
-7.07659775E-08 3.11379069E-11 2.27262660E+04 1.71124336E+01 2.47104544E+04    4
CYC5H7 Cy-1en3yl  A 9/04C  5.H  7.   0.   0.G   200.000  6000.000 1000.        1
 9.74013709E+00 2.15079576E-02-7.71169114E-06 1.24352828E-09-7.43887470E-14    2
 1.56355223E+04-2.89664925E+01 2.31203194E+00 7.01023600E-03 9.35725543E-05    3
-1.33744658E-07 5.55553794E-11 1.91721662E+04 1.72892593E+01 2.07617132E+04    4
C5H7                    C   5H   7          G    300.00   4000.00 1000.00      1        ! PREVIOUS POLIMI  CORRESPONDS TO BURCAT C5H7 Cy-1en-4-yl
 .671323690E+01 .274278890E-01-.994311090E-05 .119373240E-08 .000000000E+00    2
 .235116384E+05-.112735252E+02 .759315300E+00 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .251686000E+05 .196131100E+02                   4
RC6H9A                  C   6H   9          G    300.00   4000.00 1400.00      1
 .170842767E+02 .208842788E-01-.714529004E-05 .110943563E-08-.643676989E-13    2
 .201040204E+05-.639326012E+02-.266715213E+01 .726196475E-01-.605323920E-04    3
 .266000571E-07-.474613408E-11 .264415017E+05 .402220332E+02                   4
RCYC6H9                 C   6H   9          G    300.00   4000.00 1381.00      1
 .166730638E+02 .227088190E-01-.801509353E-05 .127088484E-08-.748275111E-13    2
 .698387216E+04-.723601536E+02-.631908086E+01 .726795534E-01-.484456826E-04    3
 .157628084E-07-.202092558E-11 .153574632E+05 .524769640E+02                   4
!HE                      HE  1               G    300.00   4000.00 1000.00      1
! .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
!-.745375000E+03 .928723974E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
! .000000000E+00 .000000000E+00-.745375000E+03 .928723974E+00                   4
HE                ATcT3EHe  1    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] He <g> ATcT ver. 1.122, DHf298 = 0.000 � 0.000 kJ/mol - fit MAR17
 2.49985609E+00 2.19365392E-07-1.07525085E-10 2.07198041E-14-1.39358612E-18    2
-7.45309155E+02 9.29535014E-01 2.49976293E+00 1.01013432E-06-8.24578465E-10    3
-6.85983306E-13 7.24751856E-16-7.45340917E+02 9.29800315E-01 0.00000000E+00    4
!AR                      AR  1               G    300.00   4000.00 1000.00      1
! .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
!-.745375000E+03 .437967491E+01 .250000000E+01 .000000000E+00 .000000000E+00    3
! .000000000E+00 .000000000E+00-.745375000E+03 .437967491E+01                   4
AR                ATcT3EAr  1    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] Ar <g> ATcT ver. 1.122, DHf298 = 0.000 � 0.000 kJ/mol - fit MAR17
 2.49989176E+00 1.56134837E-07-7.76108557E-11 1.52928085E-14-1.05304493E-18    2
-7.45328403E+02 4.38029835E+00 2.49988611E+00 2.13037960E-07 8.97320772E-10    3
-2.31395752E-12 1.30201393E-15-7.45354481E+02 4.38024367E+00 0.00000000E+00    4
!N2                      N   2               G    300.00   4000.00 1000.00      1
! .295257637E+01 .139690040E-02-.492631603E-06 .786010195E-10-.460755204E-14    2
!-.923948688E+03 .587188762E+01 .353100528E+01-.123660988E-03-.502999433E-06    3
! .243530612E-08-.140881235E-11-.104697628E+04 .296747038E+01                   4
N2                ATcT3EN   2    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] N2 <g> ATcT ver. 1.122, DHf298 = 0.000 � 0.000 kJ/mol - fit MAR17
 2.93802970E+00 1.41838030E-03-5.03281045E-07 8.07555464E-11-4.76064275E-15    2
-9.17180990E+02 5.95521985E+00 3.53603521E+00-1.58270944E-04-4.26984251E-07    3
 2.37542590E-09-1.39708206E-12-1.04749645E+03 2.94603724E+00 0.00000000E+00    4
!O2                      O   2               G    300.00   4000.00 1000.00      1
! .366096065E+01 .656365811E-03-.141149627E-06 .205797935E-10-.129913436E-14    2
!-.121597718E+04 .341536279E+01 .378245636E+01-.299673416E-02 .984730201E-05    3
!-.968129509E-08 .324372837E-11-.106394356E+04 .365767573E+01                   4
O2                ATcT3EO   2    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] O2 <g> ATcT ver. 1.122, DHf298 = 0.000 � 0.000 kJ/mol - fit MAR17
 3.65980488E+00 6.59877372E-04-1.44158172E-07 2.14656037E-11-1.36503784E-15    2
-1.21603048E+03 3.42074148E+00 3.78498258E+00-3.02002233E-03 9.92029171E-06    3
-9.77840434E-09 3.28877702E-12-1.06413589E+03 3.64780709E+00 0.00000000E+00    4
!H2                      H   2               G    300.00   4000.00  700.00      1
! .122006198E+01-.697178276E-02 .149395345E-04-.735836941E-08 .107706311E-11    2
! .964756277E+03 .127210129E+02 .000000000E+00 .000000000E+00 .000000000E+00    3
! .686975867E-08-.400441121E-11 .113556495E+04 .181719411E+02                   4
H2                ATcT3EH   2    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] H2 <g> ATcT ver. 1.122, DHf298 = 0.000 � 0.000 kJ/mol - fit MAR17
 2.90207649E+00 8.68992581E-04-1.65864430E-07 1.90851899E-11-9.31121789E-16    2
-7.97948726E+02-8.45591320E-01 2.37694204E+00 7.73916922E-03-1.88735073E-05    3
 1.95517114E-08-7.17095663E-12-9.21173081E+02 5.47184736E-01 0.00000000E+00    4
!H2O                     H   2O   1          G    300.00   4000.00 1000.00      1
! .267703890E+01 .297318160E-02-.773768890E-06 .944335140E-10-.426899910E-14    2
!-.298858940E+05 .688255000E+01 .419863520E+01-.203640170E-02 .652034160E-05    3
!-.548792690E-08 .177196800E-11-.302937260E+05-.849009010E+00                   4
H2O               ATcT3EH   2O   1    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] H2O <g> ATcT ver. 1.122, DHf298 = -241.833 � 0.027 kJ/mol - fit MAR17
 2.73117512E+00 2.95136995E-03-8.35359785E-07 1.26088593E-10-8.40531676E-15    2
-2.99169082E+04 6.55183000E+00 4.20147551E+00-2.05583546E-03 6.56547207E-06    3
-5.52906960E-09 1.78282605E-12-3.02950066E+04-8.60610906E-01-2.90858262E+04    4
!H2O2                    H   2O   2          G    300.00   4000.00 1000.00      1
! .457977305E+01 .405326003E-02-.129844730E-05 .198211400E-09-.113968792E-13    2
!-.180071775E+05 .664970694E+00 .431515149E+01-.847390622E-03 .176404323E-04    3
!-.226762944E-07 .908950158E-11-.177067437E+05 .327373319E+01                   4
H2O2              ATcT3EH   2O   2    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] H2O2 <g> ATcT ver. 1.122, DHf298 = -135.457 � 0.064 kJ/mol - fit MAR17
 4.54017480E+00 4.15970971E-03-1.30876777E-06 2.00823615E-10-1.15509243E-14    2
-1.79514029E+04 8.55881745E-01 4.23854160E+00-2.49610911E-04 1.59857901E-05    3
-2.06919945E-08 8.29766320E-12-1.76486003E+04 3.58850097E+00-1.62917334E+04    4
!CO                      C   1O   1          G    300.00   4000.00 1000.00      1
! .304848590E+01 .135172810E-02-.485794050E-06 .788536440E-10-.469807460E-14    2
!-.142661170E+05 .601709770E+01 .357953350E+01-.610353690E-03 .101681430E-05    3
! .907005860E-09-.904424490E-12-.143440860E+05 .350840930E+01                   4
CO                ATcT3EC   1O   1    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] CO <g> ATcT ver. 1.122, DHf298 = -110.523 � 0.026 kJ/mol - fit MAR17
 3.03397274E+00 1.37328118E-03-4.96445087E-07 8.10281447E-11-4.85331749E-15    2
-1.42586044E+04 6.10076092E+00 3.59508377E+00-7.21196937E-04 1.28238234E-06    3
 6.52429293E-10-8.21714806E-13-1.43448968E+04 3.44355598E+00-1.32928623E+04    4
!CO2                     C   1O   2          G    300.00   4000.00 1000.00      1
! .463651110E+01 .274145690E-02-.995897590E-06 .160386660E-09-.916198570E-14    2
!-.490249040E+05-.193489550E+01 .235681300E+01 .898412990E-02-.712206320E-05    3
! .245730080E-08-.142885480E-12-.483719710E+05 .990090350E+01                   4
CO2               ATcT3EC   1O   2    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] CO2 <g> ATcT ver. 1.122, DHf298 = -393.475 � 0.015 kJ/mol - fit MAR17
 4.63537470E+00 2.74559459E-03-9.98282389E-07 1.61013606E-10-9.22018642E-15    2
-4.90203677E+04-1.92887630E+00 2.20664321E+00 1.00970086E-02-9.96338809E-06    3
 5.47155623E-09-1.27733965E-12-4.83529864E+04 1.05261943E+01-4.73241678E+04    4
CH2O                    C   1H   2O   1     G    300.00   4000.00 1000.00      1
 .316952665E+01 .619320560E-02-.225056366E-05 .365975660E-09-.220149458E-13    2
-.145486831E+05 .604207898E+01 .479372312E+01-.990833322E-02 .373219990E-04    3
-.379285237E-07 .131772641E-10-.143791953E+05 .602798058E+00                   4
HCOOH                   C   1H   2O   2     G    300.00   4000.00 1000.00      1
 .461383160E+01 .644963640E-02-.229082510E-05 .367160470E-09-.218736750E-13    2
-.453303180E+05 .847883830E+00 .389836160E+01-.355877950E-02 .355205380E-04    3
-.438499590E-07 .171077690E-10-.467785744E+05 .734953970E+01                   4
HCO3H                   C   1H   2O   3     G    300.00   4000.00 1378.00      1
 .987503581E+01 .464663708E-02-.167230522E-05 .268624413E-09-.159595232E-13    2
-.380502456E+05-.224938942E+02 .242464726E+01 .219706380E-01-.168705546E-04    3
 .625612194E-08-.911645843E-12-.354828006E+05 .175027796E+02                   4
CH4                     C   1H   4          G    300.00   4000.00 1000.00      1
 .165326226E+01 .100263099E-01-.331661238E-05 .536483138E-09-.314696758E-13    2
-.100095936E+05 .990506283E+01 .514911468E+01-.136622009E-01 .491453921E-04    3
-.484246767E-07 .166603441E-10-.102465983E+05-.463848842E+01                   4
CH3OH                   C   1H   4O   1     G    300.00   4000.00 1000.00      1
 .352726795E+01 .103178783E-01-.362892944E-05 .577448016E-09-.342182632E-13    2
-.260028834E+05 .516758693E+01 .565851051E+01-.162983419E-01 .691938156E-04    3
-.758372926E-07 .280427550E-10-.256119736E+05-.897330508E+00                   4
CH3O2H                  C   1H   4O   2     G    300.00   4000.00 1000.00      1
 .776538058E+01 .861499712E-02-.298006935E-05 .468638071E-09-.275339255E-13    2
-.182979984E+05-.143992663E+02 .290540897E+01 .174994735E-01 .528243630E-05    3
-.252827275E-07 .134368212E-10-.168894632E+05 .113741987E+02                   4
C2H2                    C   2H   2          G    300.00   4000.00 1000.00      1
 .465878489E+01 .488396667E-02-.160828888E-05 .246974544E-09-.138605959E-13    2
 .257594042E+05-.399838194E+01 .808679682E+00 .233615762E-01-.355172234E-04    3
 .280152958E-07-.850075165E-11 .264289808E+05 .139396761E+02                   4
CH2CO                   C   2H   2O   1     G    300.00   4000.00 1000.00      1
 .575871449E+01 .635124053E-02-.225955361E-05 .362321512E-09-.215855515E-13    2
-.808533464E+04-.496490444E+01 .213241136E+01 .181319455E-01-.174093315E-04    3
 .935336040E-08-.201724844E-11-.714808520E+04 .133807969E+02                   4
CHOCHO                  C   2H   2O   2     G    300.00   4000.00 1000.00      1
 .872506895E+01 .633096819E-02-.235574814E-05 .389782853E-09-.237486912E-13    2
-.291024131E+05-.203903909E+02 .468412461E+01 .478012819E-03 .426390768E-04    3
-.579018239E-07 .231669328E-10-.271985007E+05 .451187184E+01                   4
C2H4                    C   2H   4          G    300.00   4000.00 1000.00      1
 .399182724E+01 .104833908E-01-.371721342E-05 .594628366E-09-.353630386E-13    2
 .426865851E+04-.269081762E+00 .395920063E+01-.757051373E-02 .570989993E-04    3
-.691588352E-07 .269884190E-10 .508977598E+04 .409730213E+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   4000.00 1000.00      1
 .540411080E+01 .117230590E-01-.422631370E-05 .683724510E-09-.409848630E-13    2
-.225931220E+05-.348079170E+01 .472945950E+01-.319328580E-02 .475349210E-04    3
-.574586110E-07 .219311120E-10-.215728780E+05 .410301590E+01                   4
C2H4O1-2                C   2H   4O   1     G    300.00   4000.00 1000.00      1
 .548876410E+01 .120461900E-01-.433369310E-05 .700283110E-09-.419490880E-13    2
-.918042510E+04-.707996050E+01 .375905320E+01-.944121800E-02 .803097210E-04    3
-.100807880E-06 .400399210E-10-.756081430E+04 .784974750E+01                   4
CH3CO2H                 C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .767084601E+01 .135152602E-01-.525874333E-05 .893184479E-09-.553180543E-13    2
-.557560970E+05-.154677315E+02 .278950201E+01 .999941719E-02 .342572245E-04    3
-.509031329E-07 .206222185E-10-.534752488E+05 .141053123E+02                   4
CH3OCHO                 C   2H   4O   2     G    300.00   4000.00  700.00      1
 .502910660E+01-.287377520E-01 .615808971E-04-.298073518E-07 .429774802E-11    2
-.407046731E+05 .182412180E+02 .000000000E+00 .000000000E+00 .000000000E+00    3
 .288411216E-07-.166481354E-10-.400005982E+05 .407099939E+02                   4
CH2OHCHO                C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .691088832E+01 .123280849E-01-.438373062E-05 .703055164E-09-.419009846E-13    2
-.400211587E+05-.696132551E+01 .614926095E+01-.596828114E-02 .596003337E-04    3
-.716663578E-07 .274014411E-10-.388356849E+05 .186644598E+01                   4
C2-OQOOH                C   2H   4O   3     G    300.00   4000.00 1000.00      1
 .127662941E+02 .102143437E-01-.363547001E-05 .583491588E-09-.347179974E-13    2
-.753528536E+05-.396511752E+02 .280443702E+01 .210851644E-01 .335863233E-04    3
-.702669107E-07 .326849274E-10-.720649998E+05 .151180675E+02                   4
CH3CO3H                 C   2H   4O   3     G    300.00   4000.00 1000.00      1
 .127662941E+02 .102143437E-01-.363547001E-05 .583491588E-09-.347179974E-13    2
-.753528536E+05-.396511752E+02 .280443702E+01 .210851644E-01 .335863233E-04    3
-.702669107E-07 .326849274E-10-.720649998E+05 .151180675E+02                   4
DME-OQOOH               C   2H   4O   4     G    300.00   4000.00 1000.00      1
 .114777196E+02 .831667150E-02-.185084560E-05 .103274160E-09 .000000000E+00    2
-.451075908E+05-.290204723E+02 .484746000E+01 .218580610E-01-.904284660E-05    3
 .384145300E-09 .000000000E+00-.429209100E+05 .674072600E+01                   4
C2H6                    C   2H   6          G    300.00   4000.00 1000.00      1
 .404666411E+01 .153538802E-01-.547039485E-05 .877826544E-09-.523167531E-13    2
-.124473499E+05-.968698313E+00 .429142572E+01-.550154901E-02 .599438458E-04    3
-.708466469E-07 .268685836E-10-.115222056E+05 .266678994E+01                   4
CH3OCH3                 C   2H   6O   1     G    300.00   4000.00 1000.00      1
 .564844274E+01 .163381875E-01-.586802189E-05 .946836384E-09-.566504295E-13    2
-.250864216E+05-.596267354E+01 .530562273E+01-.214253958E-02 .530873092E-04    3
-.623146897E-07 .230730916E-10-.239655820E+05 .713244569E+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   4000.00 1000.00      1
 .656243650E+01 .152042220E-01-.538967950E-05 .862250110E-09-.512897870E-13    2
-.315256210E+05-.947302020E+01 .485869570E+01-.374017260E-02 .695553780E-04    3
-.886547960E-07 .351688350E-10-.299961320E+05 .480185450E+01                   4
C2H5O2H                 C   2H   6O   2     G    300.00   4000.00 1000.00      1
 .958691079E+01 .148603589E-01-.529787964E-05 .847317148E-09-.503436325E-13    2
-.238367900E+05-.228310676E+02 .414672004E+01 .978668137E-02 .491492257E-04    3
-.742532076E-07 .311169441E-10-.214671219E+05 .984024999E+01                   4
CH2OHCH2OH              C   2H   6O   2     G    300.00   4000.00 1000.00      1
 .791471937E+01 .158415156E-01-.553486929E-05 .873346629E-09-.514003705E-13    2
-.506036554E+05-.123696999E+02 .612883088E+01-.772943096E-02 .865891028E-04    3
-.109211943E-06 .432667518E-10-.488825925E+05 .334129960E+01                   4
C3H4-P                  C   3H   4          G    300.00   4000.00 1000.00      1
 .602524000E+01 .113365420E-01-.402233910E-05 .643760630E-09-.382996350E-13    2
 .196209420E+05-.860437850E+01 .268038690E+01 .157996510E-01 .250705960E-05    3
-.136576230E-07 .661542850E-11 .208023740E+05 .987693510E+01                   4
C3H4-A                  C   3H   4          G    300.00   4000.00 1000.07      1
 .631687220E+01 .111337280E-01-.396293780E-05 .635642380E-09-.378755400E-13    2
 .201174950E+05-.109957660E+02 .261304450E+01 .121225750E-01 .185398800E-04    3
-.345251490E-07 .153350790E-10 .215415670E+05 .102261390E+02                   4
C2H3CHO                 C   3H   4O   1     G    300.00   4000.00 1000.00      1
 .820654919E+01 .128492916E-01-.464285331E-05 .751738738E-09-.451298116E-13    2
-.118838341E+05-.149881933E+02 .469868861E+01 .499965957E-02 .438587397E-04    3
-.612883900E-07 .248508985E-10-.100875286E+05 .729812046E+01                   4
CHOCH2CHO               C   3H   4O   2     G    300.00   4000.00 1000.00      1
 .104962923E+02 .120559957E-01-.434149310E-05 .699425892E-09-.418003976E-13    2
-.437332461E+05-.275425657E+02 .124227207E+01 .300698605E-01-.148206586E-05    3
-.242738150E-07 .133121686E-10-.408667843E+05 .219242842E+02                   4
CH3COCHO                C   3H   4O   2     G    300.00   4000.00 1000.00      1
 .104962923E+02 .120559957E-01-.434149310E-05 .699425892E-09-.418003976E-13    2
-.437332461E+05-.275425657E+02 .124227207E+01 .300698605E-01-.148206586E-05    3
-.242738150E-07 .133121686E-10-.408667843E+05 .219242842E+02                   4
C3H4O3                  C   3H   4O   3     G    300.00   4000.00 1388.00      1
 .137530675E+02 .108054207E-01-.364230159E-05 .560730953E-09-.323659923E-13    2
-.577839662E+05-.401019465E+02 .208981535E+01 .383715226E-01-.282590499E-04    3
 .104299134E-07-.153140407E-11-.538199819E+05 .223338530E+02                   4
KEA3BG                  C   3H   4O   4     G    300.00   4000.00 1387.00      1
 .188513241E+02 .920926912E-02-.331625639E-05 .532903065E-09-.316697392E-13    2
-.488407829E+05-.672981510E+02 .114193480E+01 .543367117E-01-.478232702E-04    3
 .206439596E-07-.352353283E-11-.431220565E+05 .263898462E+02                   4
C3H6                    C   3H   6          G    300.00   4000.00 1000.00      1
 .603870234E+01 .162963931E-01-.582130800E-05 .935936829E-09-.558603143E-13    2
-.741715057E+03-.843825992E+01 .383464468E+01 .329078952E-02 .505228001E-04    3
-.666251176E-07 .263707473E-10 .788717123E+03 .753408013E+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .811285474E+01 .171952419E-01-.606427393E-05 .967014746E-09-.573968013E-13    2
-.214419954E+05-.172623867E+02 .511393563E+01 .469115954E-02 .542574797E-04    3
-.729774751E-07 .290683409E-10-.196373114E+05 .316334698E+01                   4
C2H5CHO                 C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .744085690E+01 .177301764E-01-.634081568E-05 .102040803E-08-.609461714E-13    2
-.260055814E+05-.144195446E+02 .424529681E+01 .668296706E-02 .493337933E-04    3
-.671986124E-07 .267262347E-10-.241473007E+05 .690738560E+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .729796974E+01 .175656913E-01-.631678065E-05 .102025553E-08-.610903592E-13    2
-.295368927E+05-.127591704E+02 .555638920E+01-.283863547E-02 .705722951E-04    3
-.878130984E-07 .340290951E-10-.278325393E+05 .231960221E+01                   4
C3H6O                   C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .801491079E+01 .173919953E-01-.626027968E-05 .101188256E-08-.606239111E-13    2
-.151980838E+05-.188279964E+02 .342806676E+01 .625176642E-02 .613196311E-04    3
-.860387185E-07 .351371393E-10-.128446646E+05 .104244994E+02                   4
C3H5OOH                 C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .139268456E+02 .135384067E-01-.474335693E-05 .748389157E-09-.439105886E-13    2
-.132537727E+05-.456757848E+02 .221491505E+01 .390935107E-01-.258809564E-04    3
 .870894601E-08-.120793929E-11-.896037969E+04 .179425329E+02                   4
CH2OHCOCH3              C   3H   6O   2     G    300.00   4000.00 1000.00      1
 .110374327E+02 .169177041E-01-.598872959E-05 .957507054E-09-.569424407E-13    2
-.479270048E+05-.288076231E+02 .352624872E+01 .266034923E-01 .115090267E-04    3
-.353751170E-07 .166033210E-10-.453401970E+05 .125889401E+02                   4
CH2OHCH2CHO             C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .118936666E+02 .144153203E-01-.477525443E-05 .726036430E-09-.415285995E-13    2
-.459271652E+05-.327285750E+02 .266613285E+01 .346302298E-01-.214380719E-04    3
 .690469334E-08-.916939105E-12-.425706030E+05 .173358364E+02                   4
C3-OQOOH                C   3H   6O   3     G    300.00   4000.00 1391.00      1
 .170285271E+02 .130716784E-01-.459310856E-05 .726135156E-09-.426658337E-13    2
-.416334217E+05-.592513577E+02 .768933034E+00 .546905880E-01-.465072405E-04    3
 .203159585E-07-.358398999E-11-.363238861E+05 .268291637E+02                   4
C3H8                    C   3H   8          G    300.00   4000.00 1000.00      1
 .666919760E+01 .206108751E-01-.736512349E-05 .118434262E-08-.706914630E-13    2
-.162754066E+05-.131943379E+02 .421093013E+01 .170886504E-02 .706530164E-04    3
-.920060565E-07 .364618453E-10-.143810883E+05 .561004451E+01                   4
NC3H7OH                 C   3H   8O   1    0G   300.000  5000.000 1400.000    31 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
 1.14717073E+01 1.71812521E-02-5.78165901E-06 8.87786623E-10-5.11116063E-14    2
-3.65788256E+04-3.49774412E+01-1.28694006E-01 4.25920996E-02-2.62946409E-05    3
 8.07203568E-09-9.57756657E-13-3.24028755E+04 2.78855895E+01                   4
IC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1000.00      1
 .964183701E+01 .200230715E-01-.711967189E-05 .114138950E-08-.679935249E-13    2
-.374835623E+05-.256288343E+02 .430755345E+01 .102582798E-01 .619565411E-04    3
-.902973802E-07 .373936384E-10-.349249212E+05 .755995822E+01                   4
C3H7OOH                 C   3H   8O   2     G    300.00   4000.00 1000.00      1
 .104115631E+02 .213763889E-01-.755819870E-05 .120207180E-08-.711798090E-13    2
-.268935445E+05-.235428789E+02 .708977756E+01-.486163264E-02 .103253531E-03    3
-.133200956E-06 .530799252E-10-.244194556E+05 .174859215E+01                   4
GLYCEROL                C   3H   8O   3     G    300.00   4000.00 1000.00      1
 .143043899E+02 .198820797E-01-.705141811E-05 .112196047E-08-.663290455E-13    2
-.753417115E+05-.407500023E+02 .129036739E+01 .687295831E-01-.824160146E-04    3
 .568196772E-07-.162329302E-10-.723210175E+05 .234582202E+02                   4
!C4H2                    C   4H   2          G    300.00   4000.00 1000.00      1 !polimi
! .903147468E+01 .604725210E-02-.194878790E-05 .275486300E-09-.138560800E-13    2
! .529472934E+05-.238511290E+02 .400519100E+01 .198100000E-01-.986587660E-05    3
!-.663515820E-08 .607741290E-11 .542406400E+05 .184573600E+01                   4
C4H2                    C   4H   2          G    300.00   4000.00 1000.00      1 !Burcat kik
 8.65615648E+00 6.74465042E-03-2.36868410E-06 3.76553454E-10-2.22995205E-14    2
 5.22459295E+04-2.18462806E+01-5.02389168E-01 5.25164044E-02-9.29945578E-05    3
 8.17206506E-08-2.73537313E-11 5.38574848E+04 2.06780532E+01 5.53688672E+04    4
!C4H4                    C   4H   4          G    300.00   4000.00 1000.00      1 !ARAMCO
! .665080310E+01 .161294300E-01-.719388700E-05 .149817800E-08-.118641100E-12    2
! .311958636E+05-.979559836E+01-.191524700E+01 .527508700E-01-.716559400E-04    3
! .550724200E-07-.172862200E-10 .329785000E+05 .314199800E+02                   4
C4H4                    C   4H   4          G    300.00   4000.00 1000.00      1 !Burcat kik
 7.98456038E+00 1.20558816E-02-4.23587475E-06 6.73646140E-10-3.99059864E-14    2
 3.11993029E+04-1.67958975E+01 1.37368786E+00 2.88801256E-02-1.46863874E-05    3
-3.91045446E-09 4.78133572E-12 3.30633344E+04 1.75941274E+01 3.46213066E+04    4
FURAN                   C   4H   4O   1     G    300.00   4000.00 1000.00      1
 .135912211E+02 .987450910E-02-.345325238E-05 .544429808E-09-.319349896E-13    2
-.115639534E+05-.542513644E+02-.750030326E+01 .699899868E-01-.695485649E-04    3
 .333968809E-07-.619467883E-11-.541634292E+04 .550218432E+02                   4
CH2CCHCHO               C   4H   4O   1     G    300.00   4000.00 1000.00      1
 .929991052E+01 .152201510E-01-.615883937E-05 .112678366E-08-.769359137E-13    2
 .368009609E+04-.220663746E+02 .123852148E+01 .356054647E-01-.236786887E-04    3
 .592234361E-08 .282885884E-12 .610569242E+04 .202911558E+02                   4
C4H6  1,3-butadienT05/04C  4.H  6.   0.   0.G   200.000  6000.000 1000.        1  !Burcat MP
 7.62637466E+00 1.72523403E-02-6.09184911E-06 9.70800102E-10-5.76169721E-14    2
 9.55306395E+03-1.48325259E+01 4.10599669E+00 5.05575563E-03 5.83885454E-05    3
-8.05950198E-08 3.27447711E-11 1.15092468E+04 8.42978067E+00 1.33302095E+04    4
IC3H5CHO                C   4H   6O   1     G    300.00   4000.00 1396.00      1
 .136175682E+02 .137917192E-01-.473370118E-05 .736655226E-09-.420097974E-13    2
-.199994281E+05-.472987367E+02 .627183793E+00 .466780254E-01-.374430631E-04    3
 .158330542E-07-.273952155E-11-.157203117E+05 .216034294E+02                   4
C3H5CHO                 C   4H   6O   1     G    300.00   4000.00 1394.00      1
 .121670926E+02 .150749706E-01-.518640017E-05 .808302587E-09-.470194864E-13    2
-.156762389E+05-.365095664E+02-.227554121E-01 .441176181E-01-.322046234E-04    3
 .124986163E-07-.202269249E-11-.114618192E+05 .288193193E+02                   4
ETIBALDGB               C   4H   6O   2     G    300.00   4000.00 1000.00      1
 .130577477E+02 .906905120E-02-.308189261E-05 .476481380E-09-.275669277E-13    2
-.369274825E+05-.425273740E+02 .147485987E+00 .464706296E-01-.451901760E-04    3
 .219641008E-07-.416219125E-11-.331809255E+05 .242182934E+02                   4
ETALD4X                 C   4H   6O   2     G    300.00   4000.00 1000.00      1
 .130577477E+02 .906905120E-02-.308189261E-05 .476481380E-09-.275669277E-13    2
-.369274825E+05-.425273740E+02 .147485987E+00 .464706296E-01-.451901760E-04    3
 .219641008E-07-.416219125E-11-.331809255E+05 .242182934E+02                   4
ETIBALDGG               C   4H   6O   2     G    300.00   4000.00 1000.00      1
 .130577477E+02 .906905120E-02-.308189261E-05 .476481380E-09-.275669277E-13    2
-.369274825E+05-.425273740E+02 .147485987E+00 .464706296E-01-.451901760E-04    3
 .219641008E-07-.416219125E-11-.331809255E+05 .242182934E+02                   4
C4H6O2                  C   4H   6O   2     G    300.00   4000.00 1375.00      1
 .135393551E+02 .168328392E-01-.587873230E-05 .925553795E-09-.542254877E-13    2
-.462482008E+05-.437360830E+02 .182538964E+01 .377978336E-01-.172044878E-04    3
 .195698878E-08 .398612932E-12-.415126261E+05 .214925508E+02                   4
MACRIL                  C   4H   6O   2     G    300.00   4000.00 1000.00      1
 .962595080E+01 .202069860E-01-.684948550E-05 .109063620E-08-.671284990E-13    2
-.414857110E+05-.177414250E+02-.929250120E+00 .565245670E-01-.531143270E-04    3
 .263405850E-07-.484636380E-11-.390243280E+05 .347643170E+02                   4
KEA4X                   C   4H   6O   4     G    300.00   4000.00 1000.00      1
 .844721220E+01 .279565620E-01-.931325210E-05 .146601490E-08-.895812420E-13    2
-.149523750E+05-.219017790E+01 .170003960E+01 .665491220E-01-.743515920E-04    3
 .459831110E-07-.114108380E-10-.146870580E+05 .263355290E+02                   4
KIA4G3                  C   4H   6O   4     G    300.00   4000.00 1000.00      1
 .308381600E+02-.332377100E-02 .408622100E-05-.107259400E-08 .893684300E-13    2
-.609320200E+05-.128876900E+03 .279202700E+01 .460692000E-01-.161793100E-04    3
-.299433100E-08 .105548900E-11-.505399900E+05 .259977500E+02                   4
KIA4G2                  C   4H   6O   4     G    300.00   4000.00 1000.00      1
 .252315400E+02-.400599800E-02 .411576000E-05-.101225600E-08 .821198700E-13    2
-.541802300E+05-.106393200E+03 .276106400E+01 .360555700E-01-.139183000E-04    3
-.578268000E-09 .202447700E-12-.458617500E+05 .176080200E+02                   4
C4H8-1                  C   4H   8          G    300.00   4000.00 1392.00      1
 .113508668E+02 .180617877E-01-.616093029E-05 .954652959E-09-.553089641E-13    2
-.597871038E+04-.364369438E+02-.831372089E+00 .452580978E-01-.293658559E-04    3
 .100220436E-07-.143191680E-11-.157875035E+04 .295084236E+02                   4
IC4H8                   C   4H   8          G    300.00   4000.00 1388.00      1
 .112258330E+02 .181795798E-01-.620348592E-05 .961444458E-09-.557088057E-13    2
-.769983777E+04-.373306704E+02 .938433173E+00 .390547287E-01-.216437148E-04    3
 .587267077E-08-.614435479E-12-.374817891E+04 .191442985E+02                   4
C4H8O                   C   4H   8O   1     G    300.00   4000.00 1371.00      1
 .154228514E+02 .170211052E-01-.606347951E-05 .967354762E-09-.571992419E-13    2
-.220196123E+05-.613882135E+02-.253690104E+01 .543995707E-01-.343390305E-04    3
 .101079922E-07-.110262736E-11-.152980680E+05 .367400719E+02                   4
MEK                     C   4H   8O   1     G    300.00   4000.00 1000.00      1
 .929655016E+01 .229172746E-01-.822048591E-05 .132404838E-08-.791751980E-13    2
-.334442311E+05-.204993263E+02 .661978185E+01 .851847835E-02 .510322077E-04    3
-.658433042E-07 .249110484E-10-.315251691E+05-.109485469E+01                   4
C3H7CHO                 C   4H   8O   1     G    300.00   4000.00 1460.00      1
 .177916692E+02 .160697035E-01-.578626200E-05 .929729307E-09-.552476040E-13    2
-.343943030E+05-.708794705E+02 .269734263E+01 .347742121E-01-.145911329E-05    3
-.117722414E-07 .392653613E-11-.276350928E+05 .158339562E+02                   4
IC3H7CHO                C   4H   8O   1     G    300.00   4000.00 1391.00      1
 .137503148E+02 .183126722E-01-.628572629E-05 .978250756E-09-.568538653E-13    2
-.326938845E+05-.477281342E+02-.273021382E+00 .489696307E-01-.312770049E-04    3
 .100052945E-07-.127512074E-11-.276054737E+05 .283451139E+02                   4
!NC4H7OH                 C   4H   8O   1     G    300.00   4000.00 1000.00      1
! .863167950E+01 .241150480E-01-.832957180E-05 .134433130E-08-.835340300E-13    2
!-.230779140E+05-.163015210E+02 .173864090E+01 .369849060E-01-.680297030E-05    3
!-.128647340E-07 .662652570E-11-.209184180E+05 .207395880E+02                   4
NC4H7OH                 C   4H   8O   1     G    300.00   5000.00 1400.00      1   !Sarathy PECS c4h7oh1-1
 1.44612867E+01 1.71471992E-02-5.75989418E-06 8.83304217E-10-5.08053961E-14    2
-2.79941834E+04-5.06228722E+01-1.18168398E+00 5.97645754E-02-5.14756807E-05    3
 2.34495059E-08-4.30429836E-12-2.31416659E+04 3.12800130E+01                   4
!IC4H7OH                 C   4H   8O   1     G    300.00   4000.00 1000.00      1    !da calcolare MP
! .863167950E+01 .241150480E-01-.832957180E-05 .134433130E-08-.835340300E-13    2
!-.230779140E+05-.163015210E+02 .173864090E+01 .369849060E-01-.680297030E-05    3
!-.128647340E-07 .662652570E-11-.209184180E+05 .207395880E+02                   4
IC4H7OH                 C   4H   8O   1     G    300.00   4000.00 1384.00      1 !Sarathy PECS
 1.35043419E+01 1.78646968E-02-5.99304371E-06 9.18717641E-10-5.28435302E-14    2
-2.58255688E+04-4.44645715E+01 1.69099899E+00 4.27168891E-02-2.49281695E-05    3
 7.00961522E-09-7.23262828E-13-2.14512334E+04 1.99500833E+01                   4
ALDC6                   C   6H  12O   1     G    300.00   4000.00 1000.00      1
 .198891043E+02 .271869340E-01-.927391515E-05 .143744158E-08-.833090761E-13    2
-.397523444E+05-.760741671E+02 .137517192E+01 .665669689E-01-.404423050E-04    3
 .123836270E-07-.152905857E-11-.328740986E+05 .248343934E+02                   4
ETC3H4O2                C   3H   4O   2     G    300.00   4000.00 1404.00      1
 .130577477E+02 .906905120E-02-.308189261E-05 .476481380E-09-.275669277E-13    2
-.369274825E+05-.425273740E+02 .147485987E+00 .464706296E-01-.451901760E-04    3
 .219641008E-07-.416219125E-11-.331809255E+05 .242182934E+02                   4
RALD6XOO                C   6H  11O   3     G    300.00   3500.00 1240.00      1
 5.00092571e+01-5.34134237e-02 6.46290118e-05-2.28766994e-08 2.64030350e-12    2
-4.06673528e+04-2.20829565e+02-1.12640289e+01 1.44242337e-01-1.74470699e-04    3
 1.05671532e-07-2.32766787e-11-2.54715779e+04 8.79592018e+01                   4
RALD6X                  C   6H  11O   1     G    300.00   4000.00 1378.00      1
 1.32757019E+01	3.87287541E-02-1.48883385E-05	2.46746786E-09-1.48880472E-13    2
-1.81757665E+04-4.13894477E+01 3.91575795E+00	5.06035891E-02-1.65881567E-05    3
-1.45714100E-10	6.94235310E-13-1.35519690E+04	1.30373730E+01                   4
QA6X                    C   6H  11O   3     G    300.00   3500.00 1020.00      1
 3.16179272e+01-1.36493906e-02 3.39152683e-05-1.31900640e-08 1.56959129e-12    2
-3.26152699e+04-1.14322463e+02-3.56697724e+00 1.24330627e-01-1.68996522e-04    3
 1.19432021e-07-3.09358218e-11-2.54375494e+04 5.61211162e+01                   4
ZA6X                    C   6H  11O   5     G    300.00   3500.00 1030.00      1
 4.82844919e+01-4.15707488e-02 6.14657190e-05-2.30375151e-08 2.73823914e-12    2
-5.69207575e+04-1.98450743e+02-1.56034002e+01 2.06537570e-01-2.99857075e-04    3
 2.10828371e-07-5.40253255e-11-4.37598517e+04 1.11659856e+02                   4
KEA6X                   C   6H  10O   4     G    300.00   3500.00  890.00      1
 2.81159858e+01-1.51101039e-02 3.53666265e-05-1.35086152e-08 1.59169636e-12    2
 3.74972700e+04-9.42664402e+01 2.11579046e-01 1.10302960e-01-1.76003706e-04    3
 1.44821222e-07-4.28829769e-11 4.24642543e+04 3.71043849e+01                   4
ETALD6X                 C   6H  10O   2     G    300.00   4000.00 1000.00      1
 1.30577477E+01	9.06905120E-03-3.08189261E-06	4.76481380E-10-2.75669277E-14    2
-3.69274825E+04-4.25273740E+01 1.47485987E-01	4.64706296E-02-4.51901760E-05    3
 2.19641008E-08-4.16219125E-12-3.31809255E+04	2.42182934E+01                   4
C5H9CHO                 C   6H  10O   1     G    300.00   4000.00 1000.00      1
 .555649280E+01 .338399710E-01-.129908190E-04 .225842790E-08-.147803790E-12    2
-.155583360E+05 .376697540E+01 .117554640E+01 .506138280E-01-.305173360E-04    3
 .629100420E-08 .920183740E-12-.149438880E+05 .244076960E+02                   4
C4H7CHO                 C   6H  10O   1     G    300.00   4000.00 1000.00      1
 8.86179270E+00	2.44574708E-02-9.08860959E-06	1.53336524E-09 -9.74116382E-14   2
-1.56172875E+04-1.63712955E+01 5.76395494E-01	4.73657231E-02 -3.13609797E-05   3
 9.39481025E-09-5.51254375E-13-1.32028536E+04	2.66135077E+01                   4
HEXENOL                 C   6H  12O   1     G    300.00   4000.00 1000.00      1
 .103979970E+02 .398469010E-01-.142748760E-04 .236355490E-08-.149482190E-12    2
-.292509820E+05-.215428390E+02-.118271340E+01 .737594660E-01-.453636600E-04    3
 .102038220E-07 .738389660E-12-.264012700E+05 .372503170E+02                   4
HEXANOLOOH              C   6H  14O   3     G    300.00   4000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
RNC3OHOOX               C   3H   7O   3     G    300.00   4000.00 1000.00      1
 .411965608E+02 .371937787E-02-.401906883E-06 .401609731E-10-.217032561E-14    2
-.505341163E+05-.188000505E+03 .203813494E+01 .784218645E-01-.441306601E-04    3
 .956957259E-08-.134730026E-11-.362640104E+05 .268180208E+02                   4
QNC3OHOOX               C   3H   7O   3     G    300.00   4000.00 1000.00      1
 .410726584E+02 .325163393E-02-.312770829E-06 .282397537E-10-.137453673E-14    2
-.449667530E+05-.183380687E+03 .255294420E+01 .839412693E-01-.653740910E-04    3
 .319006074E-07-.896548855E-11-.312800193E+05 .261620056E+02                   4
ZNC3OHOOX               C   3H   7O   5     G    300.00   4000.00 1000.00      1
 .164918847E+02 .468250506E-01-.164871837E-04 .270739186E-08-.170379572E-12    2
-.513214862E+05-.386393956E+02 .131429341E+01 .103179790E+00-.802039006E-04    3
 .264187232E-07-.137184908E-11-.487698967E+05 .341039048E+02                   4
KEHYNC3OH               C   3H   6O   4     G    300.00   4000.00 1000.00      1
 .603831357E+00 .666768020E-01-.271765190E-04 .493142950E-08-.332781746E-12    2
-.637785333E+05 .469431419E+02 .227567354E+01 .864199139E-01-.619813992E-04    3
 .165976198E-07 .130342673E-11-.669640942E+05 .287560117E+02                   4
KEA3B3L                 C   3H   4O   4     G    300.00   4000.00 1387.00      1
 .188513241E+02 .920926912E-02-.331625639E-05 .532903065E-09-.316697392E-13    2
-.488407829E+05-.672981510E+02 .114193480E+01 .543367117E-01-.478232702E-04    3
 .206439596E-07-.352353283E-11-.431220565E+05 .263898462E+02                   4
!************************Hexanol Thermo*********************************!         !MP
C6H13OH                 C   6H  14O   1     G    300.00   4000.00 1000.00      1
 .215498620E+02 .270477890E-01-.794877720E-05 .114579960E-08-.659841990E-13    2
-.486288910E+05-.832675700E+02 .811415610E+00 .696693440E-01-.335770780E-04    3
 .354337360E-08 .127138890E-11-.415253200E+05 .290476130E+02                   4
RHEX1OHA                C   6H  13O   1     G    300.00   4000.00 1000.00      1
 .224822920E+02 .220633650E-01-.560837910E-05 .726127710E-09-.387814070E-13    2
-.271730000E+05-.857930980E+02 .712225620E+00 .741183910E-01-.546395530E-04    3
 .255721450E-07-.612147960E-11-.200816860E+05 .302884250E+02                   4
RHEX1OHB                C   6H  13O   1     G    300.00   4000.00 1000.00      1
 .226977810E+02 .216816440E-01-.545814460E-05 .701621370E-09-.372876710E-13    2
-.252458440E+05-.868857500E+02-.372279850E+00 .818340110E-01-.718173030E-04    3
 .412142000E-07-.112622190E-10-.180154040E+05 .348058320E+02                   4
RESAN1OHC               C   6H  13O   1     G    300.00   4000.00 1000.00      1
 .226977810E+02 .216816440E-01-.545814460E-05 .701621370E-09-.372876710E-13    2
-.252458440E+05-.868857500E+02-.372279850E+00 .818340110E-01-.718173030E-04    3
 .412142000E-07-.112622190E-10-.180154040E+05 .348058320E+02                   4
RESAN1OHD               C   6H  13O   1     G    300.00   4000.00 1000.00      1
 .226977810E+02 .216816440E-01-.545814460E-05 .701621370E-09-.372876710E-13    2
-.252458440E+05-.868857500E+02-.372279850E+00 .818340110E-01-.718173030E-04    3
 .412142000E-07-.112622190E-10-.180154040E+05 .348058320E+02                   4
RESAN1OHE               C   6H  13O   1     G    300.00   4000.00 1000.00      1
 .224920710E+02 .220734010E-01-.562121570E-05 .729891430E-09-.391193430E-13    2
-.252098520E+05-.858406450E+02 .712452890E+00 .741594210E-01-.545500620E-04    3
 .253264660E-07-.599609950E-11-.181213770E+05 .302764260E+02                   4
RESAN1OHF               C   6H  13O   1     G    300.00   4000.00 1000.00      1
 .230495220E+02 .216574500E-01-.550175860E-05 .714146520E-09-.383251170E-13    2
-.243130620E+05-.891266780E+02-.208731200E+00 .797328870E-01-.641229850E-04    3
 .327538710E-07-.826671460E-11-.169163750E+05 .341480100E+02                   4
RESAN1O                 C   6H  13O   1     G    300.00   4000.00 1000.00      1
 .223293590E+02 .231753250E-01-.612610670E-05 .818680350E-09-.448138400E-13    2
-.230509100E+05-.883801270E+02-.599555790E+00 .741732340E-01-.454306210E-04    3
 .140138330E-07-.200701590E-11-.154257910E+05 .347537120E+02                   4
!
QC6OHOOX                C   6H  13O   3     G    300.00   4000.00 1000.00      1
 .410726584E+02 .325163393E-02-.312770829E-06 .282397537E-10-.137453673E-14    2
-.449667530E+05-.183380687E+03 .255294420E+01 .839412693E-01-.653740910E-04    3
 .319006074E-07-.896548855E-11-.312800193E+05 .261620056E+02                   4
RC6OHOOX                C   6H  13O   3     G    300.00   4000.00 1000.00      1
 .411965608E+02 .371937787E-02-.401906883E-06 .401609731E-10-.217032561E-14    2
-.505341163E+05-.188000505E+03 .203813494E+01 .784218645E-01-.441306601E-04    3
 .956957259E-08-.134730026E-11-.362640104E+05 .268180208E+02                   4
ZC6OHOOX                C   6H  13O   5     G    300.00   4000.00 1000.00      1
 .164918847E+02 .468250506E-01-.164871837E-04 .270739186E-08-.170379572E-12    2
-.513214862E+05-.386393956E+02 .131429341E+01 .103179790E+00-.802039006E-04    3
 .264187232E-07-.137184908E-11-.487698967E+05 .341039048E+02                   4
ETALD6                  C   6H  12O   2     G    300.00   4000.00 1393.00      1
 .134576640E+02 .361254510E-01-.126982530E-04 .207621190E-08-.130253340E-12    2
-.276938870E+05-.443481370E+02-.480166100E+01 .824119080E-01-.502893530E-04    3
 .107391800E-07 .748536430E-12-.223889220E+05 .511845550E+02                   4
KEHYC6OH                C   6H  12O   4     G    300.00   4000.00 1000.00      1
 .603831357E+00 .666768020E-01-.271765190E-04 .493142950E-08-.332781746E-12    2
-.637785333E+05 .469431419E+02 .227567354E+01 .864199139E-01-.619813992E-04    3
 .165976198E-07 .130342673E-11-.669640942E+05 .287560117E+02                   4
! 
NC4-OQOOH               C   4H   8O   3     G    300.00   4000.00 1388.00      1
 .195955254E+02 .180568312E-01-.629994700E-05 .991157547E-09-.580382406E-13    2
-.461054913E+05-.709333761E+02 .243440296E+01 .605409309E-01-.481250984E-04    3
 .203656751E-07-.357059537E-11-.402872220E+05 .205488821E+02                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   4000.00 1390.00      1
 .195047991E+02 .181701803E-01-.634838146E-05 .999797067E-09-.585883751E-13    2
-.450007951E+05-.705122130E+02 .549934041E+00 .642751153E-01-.501779820E-04    3
 .203546231E-07-.338767418E-11-.385647626E+05 .307013051E+02                   4
KEHYBU1                 C   4H   8O   4     G    300.00   4000.00 1396.00      1
 .219367270E+02 .180406285E-01-.626171080E-05 .981855896E-09-.573639516E-13    2
-.664546784E+05-.813588272E+02-.445736457E+01 .947202096E-01-.937478682E-04    3
 .464802131E-07-.899314409E-11-.587131282E+05 .551970961E+02                   4
IC4H10                  C   4H  10          G    300.00   4000.00 1000.00      1
 .508434390E+01 .331851280E-01-.124047670E-04 .152753620E-08 .000000000E+00    2
-.195243797E+05-.392308050E+01-.128398800E+01 .519486400E-01-.308267920E-04    3
 .755438110E-08 .000000000E+00-.179038400E+05 .285063500E+02                   4
!NC4H10                  C   4H  10          G    300.00   4000.00 1000.00      1
NC4H10                  C   4H  10          G    300.00   4000.00 1000.00      1
 .105251152E+02 .235908740E-01-.785389060E-05 .114561140E-08-.599309560E-13    2
-.204952316E+05-.321928008E+02 .157641510E+01 .345897230E-01 .697016090E-05    3
-.281636370E-07 .123751170E-10-.171470040E+05 .178727420E+02                   4
N1C4H9OH                C   4H  10O   1     G   300.000  5000.000 1400.000     1 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 12_08_2016_14_12_47
+1.48022849E+01+2.15268606E-02-7.27127618E-06+1.11937370E-09-6.45600513E-14    2
-4.07592510E+04-5.13528547E+01-4.59550266E-01+5.55978022E-02-3.56641050E-05    3
+1.15878847E-08-1.49962538E-12-3.53225632E+04+3.11360441E+01+0.00000000E+00    4
N2C4H9OH                C   4H  10O   1     G    300.00   4000.00 1390.00      1
 .151582366E+02 .215048627E-01-.741631184E-05 .115764678E-08-.674130532E-13    2
-.429113728E+05-.549620416E+02-.304705097E+00 .567446943E-01-.387293873E-04    3
 .141775813E-07-.220696859E-11-.373601662E+05 .285520284E+02                   4
TC4H9OH                 C   4H  10O   1     G    300.00   4000.00 1395.00      1
 .151183592E+02 .214941230E-01-.730928419E-05 .113021881E-08-.653833962E-13    2
-.450124898E+05-.575375902E+02-.861795957E+00 .603867730E-01-.445191256E-04    3
 .177406426E-07-.295852901E-11-.395611057E+05 .278278048E+02                   4
IC4H9OH                 C   4H  10O   1     G    300.00   4000.00 1426.00      1
 .145203606E+02 .218826590E-01-.741886985E-05 .114493281E-08-.661481541E-13    2
-.415815847E+05-.516504190E+02-.808654483E+00 .568695746E-01-.379891888E-04    3
 .133635469E-07-.195588405E-11-.361485459E+05 .310126347E+02                   4
C4H9OOH                 C   4H  10O   2     G    300.00   4000.00 1389.00      1
 .182257559E+02 .215996217E-01-.748424942E-05 .117205153E-08-.684096331E-13    2
-.342341151E+05-.670536388E+02 .607792497E+00 .624669916E-01-.444490375E-04    3
 .167754668E-07-.265938189E-11-.280070327E+05 .278025473E+02                   4
C5H4O Cy CPD-ONE  T 3/10C  5.H  4.O  1.   0.G   200.000  6000.000 1000.        1  !C3 MECH
 1.00806850E+01 1.61143434E-02-5.83314395E-06 9.46759172E-10-5.68972158E-14    2     
 1.94364640E+03-2.94552495E+01 2.64575563E-01 3.34873926E-02 1.67735280E-06    3
-2.96207072E-08 1.54431326E-11 5.11159292E+03 2.35378826E+01 6.64245999E+03    4
!CYC5H4O                 C   5H   4O   1     G    300.00   4000.00 1000.00      1   ! DH similar to C5H4O new at low T, but bery different Cp
! .558734350E+01 .254149730E-01-.929145880E-05 .112347330E-08 .000000000E+00    2
! .339172461E+04-.552979995E+01-.427809100E+01 .546170700E-01-.380993520E-04    3
! .105947040E-07 .000000000E+00 .589093400E+04 .446629800E+02                   4
! YOMMEE JPCA 120 (2016) 433-451
C5H3O-3           ---LITH   3O   1C   5     G     300.0    5000.0  1401.0      1
   1.29591933E1  1.02293393E-2 -3.53287746E-6 5.52201896E-10-3.21926864E-14    2
   3.17665892E4  -4.38962623E1  -2.04669181E0  5.20908055E-2 -4.90700703E-5    3
  2.31483526E-8-4.28871558E-12   3.62791216E4   3.42501989E1                   4
FURFURAL                C   5H   4O   2     G    300.00   4000.00 1000.00      1
 .159553578E+02 .122096134E-01-.419491662E-05 .654219009E-09-.381060338E-13    2
-.255664634E+05-.596830465E+02-.186260023E+01 .570946426E-01-.476338594E-04    3
 .197949337E-07-.326585828E-11-.197873020E+05 .347179869E+02                   4
CYC5H6                  C   5H   6          G    300.00   4000.00 1000.00      1
 .230537462E+00 .409571826E-01-.241588958E-04 .679763480E-08-.736374421E-12    2
 .143779465E+05 .202551234E+02-.513691194E+01 .606953453E-01-.460552837E-04    3
 .128457201E-07 .741214852E-12 .153675713E+05 .461567559E+02                   4
MEFU2                   C   5H   6O   1     G    300.00   4000.00 1000.00      1
 .459933100E+01 .340025700E-01-.175181400E-04 .423464670E-08-.375757330E-12    2
-.129526080E+05 .466753790E+00-.284971730E+01 .552316440E-01-.365110720E-04    3
 .832948240E-08 .742313490E-12-.110344430E+05 .385458850E+02                   4
C5H8                    C   5H   8          G    300.00   4000.00 1000.00      1
 .797205310E+01 .268614160E-01-.956546320E-05 .113079120E-08 .000000000E+00    2
 .510466811E+04-.185090870E+02 .176636500E+01 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .684030700E+04 .137180600E+02                   4
CYC5H8                  C   5H   8          G    300.00   4000.00 1000.00      1
 .772447728E+01 .283223160E-01-.115452360E-04 .215408150E-08-.150541780E-12    2
-.782614232E+03-.197696844E+02 .268981400E+01 .209545500E-02 .113036870E-03    3
-.154080700E-06 .627636580E-10 .231396630E+04 .152940560E+02                   4
C5H8O                   C   5H   8O   1     G    300.00   4000.00 1000.00      1
 .154011002E+02 .203490440E-01-.699742510E-05 .109031908E-08-.634192782E-13    2
-.910076428E+04-.580710041E+02-.514624016E+01 .722177875E-01-.580157542E-04    3
 .242093068E-07-.410120178E-11-.236133441E+04 .508920452E+02                   4
MCROT                   C   5H   8O   2     G    300.00   4000.00 1000.00      1
 .110840220E+02 .266681570E-01-.910298150E-05 .145819250E-08-.902072000E-13    2
-.461868520E+05-.238654710E+02 .115411390E+01 .550597160E-01-.356332020E-04    3
 .867407750E-08 .746845670E-12-.435806950E+05 .269868980E+02                   4
ETMB583                 C   5H   8O   3     G    300.00   4000.00 1000.00      1
 .164044820E+02 .257082970E-01-.901921340E-05 .147114070E-08-.920586850E-13    2
-.622657890E+05-.550660710E+02-.249091940E+01 .790685040E-01-.564648800E-04    3
 .115540360E-07 .278656790E-11-.573317190E+05 .417407460E+02                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   4000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5H8O4                  C   5H   8O   4     G    300.00   4000.00 1000.00      1
 .217298154E+02 .217807665E-01-.749545594E-05 .116860895E-08-.680038942E-13    2
-.866505360E+05-.835752527E+02-.684199090E+01 .100610553E+00-.924172541E-04    3
 .429800586E-07-.789719358E-11-.779623201E+05 .655426910E+02                   4
KEHYMB                  C   5H   8O   5     G    300.00   4000.00 1000.00      1
 .130410150E+02 .302430520E-01-.103682550E-04 .166520830E-08-.103159200E-12    2
-.605793360E+05-.352927630E+02-.187604440E+01 .779613480E-01-.656695630E-04    3
 .280818550E-07-.405575270E-11-.569013010E+05 .398655930E+02                   4
B1M3                    C   5H  10          G    300.00   4000.00 1394.00      1
 .144242929E+02 .226454984E-01-.773646334E-05 .119999861E-08-.695711276E-13    2
-.114981027E+05-.530391197E+02-.964397004E+00 .568482691E-01-.366324275E-04    3
 .123008921E-07-.171392531E-11-.593502026E+04 .302998433E+02                   4
B2M2                    C   5H  10          G    300.00   4000.00 1389.00      1
 .140426423E+02 .227915348E-01-.774902598E-05 .119814522E-08-.693127003E-13    2
-.132160483E+05-.514469569E+02 .604882839E+00 .496635256E-01-.266571142E-04    3
 .647312078E-08-.484017883E-12-.806312207E+04 .223818263E+02                   4
B1M2                    C   5H  10          G    300.00   4000.00 1392.00      1
 .141931279E+02 .226551019E-01-.770008627E-05 .119031326E-08-.688489604E-13    2
-.119491010E+05-.510688681E+02-.539429136E+00 .544489715E-01-.332707895E-04    3
 .103047694E-07-.128363329E-11-.653967251E+04 .290349986E+02                   4
NC5H10                  C   5H  10          G    300.00   4000.00 1389.00      1
 .141108203E+02 .228348272E-01-.778626835E-05 .120627491E-08-.698795983E-13    2
-.114335029E+05-.501593461E+02-.541560551E+00 .539629918E-01-.323508738E-04    3
 .977416037E-08-.118534668E-11-.598606169E+04 .297142748E+02                   4
C4H9CHO                 C   5H  10O   1     G    300.00   4000.00 1507.00      1
 .197928063E+02 .217870723E-01-.780397879E-05 .124956209E-08-.740724001E-13    2
-.382553694E+05-.801632581E+02 .392970436E+01 .374486092E-01 .427678157E-05    3
-.168019085E-07 .508443447E-11-.306588984E+05 .125431056E+02                   4
RALD5X                  C   5H   9O   1     G    300.00   4000.00 1517.00      1   
 .190577032E+02 .197405268E-01-.706907553E-05 .113169306E-08-.670771090E-13    2
-.128899482E+05-.729817022E+02 .467212037E+01 .343554368E-01 .295219352E-05    3
-.145463894E-07 .444316435E-11-.603466621E+04 .109564879E+02                   4 
RALD5XOO                C   5H   9O   3     G    300.00   3500.00 1240.00      1   
 5.00092571e+01-5.34134237e-02 6.46290118e-05-2.28766994e-08 2.64030350e-12    2
-4.06673528e+04-2.20829565e+02-1.12640289e+01 1.44242337e-01-1.74470699e-04    3
 1.05671532e-07-2.32766787e-11-2.54715779e+04 8.79592018e+01                   4
RALD5X                  C   5H   9O   1     G    300.00   4000.00 1378.00      1   
 1.32757019E+01	3.87287541E-02-1.48883385E-05	2.46746786E-09-1.48880472E-13    2
-1.81757665E+04-4.13894477E+01 3.91575795E+00	5.06035891E-02-1.65881567E-05    3
-1.45714100E-10	6.94235310E-13-1.35519690E+04	1.30373730E+01                   4
QA5X                    C   5H   9O   3     G    300.00   3500.00 1020.00      1   
 3.16179272e+01-1.36493906e-02 3.39152683e-05-1.31900640e-08 1.56959129e-12    2
-3.26152699e+04-1.14322463e+02-3.56697724e+00 1.24330627e-01-1.68996522e-04    3
 1.19432021e-07-3.09358218e-11-2.54375494e+04 5.61211162e+01                   4
ZA5X                    C   5H   9O   5     G    300.00   3500.00 1030.00      1   
 4.82844919e+01-4.15707488e-02 6.14657190e-05-2.30375151e-08 2.73823914e-12    2
-5.69207575e+04-1.98450743e+02-1.56034002e+01 2.06537570e-01-2.99857075e-04    3
 2.10828371e-07-5.40253255e-11-4.37598517e+04 1.11659856e+02                   4
KEA5X                   C   5H   8O   4     G    300.00   3500.00  890.00      1   
 2.81159858e+01-1.51101039e-02 3.53666265e-05-1.35086152e-08 1.59169636e-12    2
 3.74972700e+04-9.42664402e+01 2.11579046e-01 1.10302960e-01-1.76003706e-04    3
 1.44821222e-07-4.28829769e-11 4.24642543e+04 3.71043849e+01                   4
IC4H9CHO                C   5H  10O   1     G    300.00   4000.00 1383.00      1
 .170194059E+02 .223541546E-01-.759760895E-05 .117496754E-08-.679975164E-13    2
-.369143302E+05-.635871575E+02 .861033163E+00 .573441683E-01-.359178644E-04    3
 .113951893E-07-.146205706E-11-.309951354E+05 .242264151E+02                   4
!C5H9OH                  C   5H  10O   1     G    300.00   4000.00 1000.00      1
! .107143420E+02 .300909990E-01-.104241840E-04 .168678680E-08-.105053190E-12    2
!-.266832230E+05-.257609100E+02-.581915140E+00 .590151210E-01-.307994630E-04    3
! .522248800E-09 .379832970E-11-.235468110E+05 .329467200E+02                   4
C5H9OH                  C   5H  10O   1     G    300.00   5000.00 1404.00      1 !Sarahty pecs 2015, c5h9oh1-1
 1.88402399E+01 2.07213749E-02-7.00668162E-06 1.07917426E-09-6.22553029E-14    2
-3.24792357E+04-7.37908378E+01-3.75711664E+00 8.61350068E-02-8.11095643E-05    3
 3.92658441E-08-7.48846199E-12-2.58553432E+04 4.31553562E+01                   4
!IC5H9OH                 C   5H  10O   1     G    300.00   4000.00 1394.00      1
! .147423131E+02 .219843767E-01-.751584192E-05 .116633393E-08-.676421638E-13    2
!-.416616600E+05-.528466211E+02-.837465362E+00 .576520639E-01-.390215462E-04    3
! .140131231E-07-.211159111E-11-.361265628E+05 .311701525E+02                   4
IC5H9OH                 C   5H  10O   1     G    300.00   5000.00 1401.00      1 !Sarahty pecs 2015, ic5h9oh1-1
 1.72230301E+01 2.22593435E-02-7.57391529E-06 1.17156666E-09-6.77917454E-14    2
-3.31186152E+04-6.50020716E+01-1.94022087E+00 7.14827733E-02-5.72564918E-05    3
 2.43814756E-08-4.24851023E-12-2.68798428E+04 3.63828341E+01                   4
NC5H10-O                C   5H  10O   1     G    300.00   4000.00 1373.00      1
 .187152768E+02 .216122625E-01-.768638433E-05 .122492227E-08-.723734176E-13    2
-.274341627E+05-.786690289E+02-.351633623E+01 .686975884E-01-.446579237E-04    3
 .140670556E-07-.174934766E-11-.191663581E+05 .425589840E+02                   4
NEOC5H10-O              C   5H  10O   1     G    300.00   4000.00 1406.00      1
 .182053093E+02 .222888126E-01-.759419141E-05 .117633164E-08-.681511068E-13    2
-.260973639E+05-.785614741E+02-.704702259E+01 .864172552E-01-.702610933E-04    3
 .290540959E-07-.480586102E-11-.179483330E+05 .550571499E+02                   4
CH3OCH3                 C   2H   6O   1    0G    300.00   5000.00 1999.00      1!21 U. Burke
 6.03232751e+00 1.56155270e-02-5.50761030e-06 8.75666140e-10-5.17180562e-14    2
-2.52690354e+04-8.25885183e+00 2.05597390e+00 2.07019456e-02-5.00382376e-06    3
-1.62279885e-09 6.84330155e-13-2.35494445e+04 1.45029944e+01                   4 
CH3OCH2                 C   2H   5O   1    0G    300.00   5000.00 1395.00      1!11  U. Burke
 6.62621974e+00 1.22219496e-02-4.12416696e-06 6.34127512e-10-3.65317390e-14    2
-3.33965890e+03-8.95305753e+00 1.58874948e+00 2.24414123e-02-1.19434933e-05    3
 3.37160213e-09-4.15077249e-13-1.37208255e+03 1.87548958e+01                   4
DME-OO                  C   2H   5O   3    0G    300.00  5000.00 1441.00       1!21  U. Burke
 1.19179361e+01 1.19412867e-02-3.93526185e-06 5.95756132e-10-3.39597705e-14    2
-2.34231833e+04-3.20096863e+01 3.39930541e+00 3.09460407e-02-1.92548181e-05    3
 5.76033887e-09-6.16081571e-13-2.04433218e+04 1.39429608e+01                   4
DME-QOOH                C   2H   5O   3    0G    300.00  5000.00 1418.00       1!21 U. Burke
 1.23892901e+01 1.11758961e-02-3.59249095e-06 5.34196366e-10-3.00536541e-14    2
-1.80551598e+04-3.29576862e+01 1.62245477e-01 4.76101093e-02-4.52046954e-05    3
 2.18379311e-08-4.11295947e-12-1.46498100e+04 2.98253164e+01                   4
DME-OOQOOH              C   2H   5O   5    0G    300.00  5000.00 1433.00       1!31 U. Burke
 1.77378326e+01 1.13589899e-02-3.67382539e-06 5.49255712e-10-3.10405899e-14    2
-3.82903058e+04-5.66609932e+01 2.39977678e+00 5.39881943e-02-4.87969524e-05    3
 2.19792134e-08-3.86106979e-12-3.37824638e+04 2.30683371e+01                   4
DME-OQOOH               C   2H   4O   4    0G    300.00  5000.00  1386.00      1!31 U. Burke
 1.57136128e+01 9.64430166e-03-3.44136025e-06 5.49722196e-10-3.25360322e-14    2
-6.29409094e+04-5.29505242e+01 1.21909586e+00 4.28858235e-02-3.17634222e-05    3
 1.11542676e-08-1.49753153e-12-5.79287926e+04 2.49759193e+01                   4
MTBE-O                  C   5H  10O   2     G    300.00   4000.00 1397.00      1
 .193844587E+02 .224929046E-01-.748169734E-05 .114123661E-08-.654437288E-13    2
-.558416627E+05-.795832532E+02-.518049059E+01 .839546669E-01-.663790553E-04    3
 .267623941E-07-.432034827E-11-.478415885E+05 .506953652E+02                   4
MB                      C   5H  10O   2     G    300.00   4000.00 1380.00      1
 .190094725E+02 .236503722E-01-.822978452E-05 .129246265E-08-.755862836E-13    2
-.634989152E+05-.732469099E+02 .316208825E+01 .552915358E-01-.311610102E-04    3
 .842394129E-08-.872222021E-12-.573385240E+05 .139723817E+02                   4
NEOC5-OQOOH             C   5H  10O   3     G    300.00   4000.00 1397.00      1
 .237028187E+02 .215843890E-01-.747470111E-05 .117038715E-08-.683143724E-13    2
-.509464263E+05-.948314143E+02 .101097520E+01 .753376897E-01-.559848192E-04    3
 .210040666E-07-.316727025E-11-.432003697E+05 .266737910E+02                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   4000.00 1389.00      1
 .227422860E+02 .225948063E-01-.786379640E-05 .123514506E-08-.722413862E-13    2
-.501979972E+05-.864068664E+02 .227305950E+01 .724929431E-01-.560597536E-04    3
 .231254746E-07-.397203084E-11-.431866364E+05 .229745558E+02                   4
MTBE-OQOOH              C   5H  10O   4     G    300.00   4000.00 1386.00      1
 .259492704E+02 .217762181E-01-.754080079E-05 .118109778E-08-.689663912E-13    2
-.659884236E+05-.102260628E+03 .215705064E+01 .770950997E-01-.562944956E-04    3
 .205751475E-07-.301215733E-11-.577585957E+05 .255153989E+02                   4
KEHYP1OH                C   5H  10O   4     G    300.00   4000.00 1391.00      1
 .241671480E+02 .230357774E-01-.791201902E-05 .123189743E-08-.716178065E-13    2
-.696422759E+05-.907717133E+02 .209051128E+01 .771281020E-01-.592331258E-04    3
 .236078672E-07-.383619864E-11-.622442740E+05 .268708461E+02                   4
KEHYIPOH                C   5H  10O   4     G    300.00   4000.00 1391.00      1
 .254040364E+02 .213220358E-01-.718760689E-05 .110596704E-08-.637962798E-13    2
-.743944256E+05-.957197841E+02 .249561727E+01 .809896491E-01-.680713112E-04    3
 .297755952E-07-.525877030E-11-.670549235E+05 .251315082E+02                   4
NC5H12                  C   5H  12          G    300.00   4000.00 1000.00      1
 .142233709E+02 .264253600E-01-.834599270E-05 .125651470E-08-.740004510E-13    2
-.247106388E+05-.503994927E+02-.393634560E+00 .578781330E-01-.285392090E-04    3
 .347472500E-08 .106523800E-11-.198713480E+05 .281908260E+02                   4
NEOC5H12                C   5H  12          G    300.00   4000.00 1397.00      1
 .174488013E+02 .245462377E-01-.835182479E-05 .129219708E-08-.747942850E-13    2
-.292378530E+05-.754164601E+02-.288372771E+01 .722417687E-01-.511106166E-04    3
 .187342407E-07-.280628313E-11-.222171069E+05 .336765462E+02                   4
MTBE                    C   5H  12O   1     G    300.00   4000.00 1000.00      1
 .888656643E+01 .420057870E-01-.178904220E-04 .345077750E-08-.247674430E-12    2
-.405353691E+05-.208281992E+02-.162610860E+01 .742240170E-01-.539682020E-04    3
 .210023490E-07-.342702090E-11-.378579060E+05 .325557600E+02                   4
IC5H11OH                C   5H  12O   1     G    300.00   4000.00 1394.00      1
 .176659926E+02 .264001578E-01-.897091677E-05 .138657980E-08-.801947316E-13    2
-.458703080E+05-.669958017E+02-.997731650E+00 .689216907E-01-.460606099E-04    3
 .161906169E-07-.236803054E-11-.392443688E+05 .336827033E+02                   4
C5H11OH                 C   5H  12O   1    0G   300.000  5000.000 1399.000    51 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
 1.81326422E+01 2.58734469E-02-8.76147510E-06 1.35108218E-09-7.80169568E-14    2
-4.49393846E+04-6.77258765E+01-7.40082990E-01 6.83880275E-02-4.47177434E-05    3
 1.49115071E-08-1.99981896E-12-3.82501077E+04 3.41515985E+01                   4
NC5H11OOH               C   5H  12O   2     G    300.00   4000.00 1391.00      1
 .215962451E+02 .259122865E-01-.896302814E-05 .140202940E-08-.817685827E-13    2
-.395542326E+05-.852046644E+02-.443227141E+00 .781363104E-01-.573273118E-04    3
 .222802059E-07-.361215684E-11-.318952281E+05 .330316890E+02                   4
!C6H2                    C   6H   2          G    300.00   4000.00 1000.00      1 !polimi
! .127565190E+02 .803438100E-02-.261821500E-05 .372506000E-09-.187885000E-13    2
! .807546900E+05-.404126200E+02 .575108500E+01 .263671900E-01-.116675960E-04    3
!-.107144980E-07 .879029700E-11 .826201200E+05-.433553200E+01                   4
C6H2              T 8/10C   6H   2    0    0G   200.000  6000.000 1000.        1 !Burcat kik
 1.25237986E+01 8.78597449E-03-3.13663802E-06 5.04347263E-10-3.01110703E-14    2
 7.97838798E+04-3.88501187E+01-5.94408010E-01 7.46613698E-02-1.35848115E-04    3
 1.22198283E-07-4.17697584E-11 8.21259933E+04 2.21178523E+01 8.42887915E+04    4
!BENZYNE                 C   6H   4          G    300.00   4000.00 1000.00      1 !polimi
! .105707063E+02 .156860613E-01-.568267148E-05 .922956737E-09-.554966417E-13    2
! .504976657E+05-.332563927E+02 .721604591E+00 .247976151E-01 .316372209E-04    3
!-.653230986E-07 .296082142E-10 .539797980E+05 .216733825E+02                   4
CYC6H4                  C   6H   4          G    300.00   4000.00 1000.00      1 !Burcat kik
 1.05707063E+01 1.56860613E-02-5.68267148E-06 9.22956737E-10-5.54966417E-14    2
 5.04976657E+04-3.32563927E+01 7.21604591E-01 2.47976151E-02 3.16372209E-05    3
-6.53230986E-08 2.96082142E-11 5.39797980E+04 2.16733825E+01 5.54615216E+04    4
LC6H4                   C   6H   4          G    300.00   4000.00 1000.00      1
 .171831170E+02 .664876580E-02-.124162630E-05 .146974480E-09-.913980130E-14    2
 .550769540E+05-.644351830E+02 .193231390E+01 .390321830E-01-.692271090E-05    3
-.270933570E-07 .157302520E-10 .596919480E+05 .165160230E+02                   4
O-C6H4O2                H  4 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! DHof -16.68 LPM automech from C6H5+O2 paper
 8.42783350E+00 3.06980473E-02-1.61682962E-05 4.08466242E-09-4.02066090E-13    2
-1.43573182E+04-1.83737356E+01 9.58195510E-01 4.14373472E-02 3.16843114E-06    3
-3.90359010E-08 2.01121081E-11-1.20255999E+04 2.20620096E+01                   4
C6H4O2                  H  4 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! DHof -24.55 LPM automech from C6H5+O2 paper
 8.46782730E+00 3.06456600E-02-1.61417824E-05 4.07864825E-09-4.01557746E-13    2
-1.83291516E+04-1.94722053E+01 9.59943977E-01 4.15600573E-02 2.96367471E-06    3
-3.89598489E-08 2.01249683E-11-1.59926336E+04 2.11378236E+01                   4
!C6H6                    C   6H   6          G    300.00   4000.00 1000.00      1 !polimi 
! .129109067E+02 .172329600E-01-.502421020E-05 .589349680E-09-.194752100E-13    2
! .366437279E+04-.500281184E+02-.313801200E+01 .472310300E-01-.296220700E-05    3
!-.326281900E-07 .171869100E-10 .889003000E+04 .365757300E+02                   4
C6H6                    C   6H   6          G    300.00   4000.00 1000.00      1! Burcat kik
 1.10809576E+01 2.07176746E-02-7.52145991E-06 1.22320984E-09-7.36091279E-14    2
 4.30641035E+03-4.00413310E+01 5.04818632E-01 1.85020642E-02 7.38345881E-05    3
-1.18135741E-07 5.07210429E-11 8.55247913E+03 2.16412893E+01 9.96811598E+03    4
LC6H6                   C   6H   6          G    300.00   4000.00 1000.00      1
 .133755312E+02 .181053970E-01-.671790940E-05 .114930710E-08-.753903640E-13    2
 .353349989E+05-.436278915E+02-.284372350E+01 .754240600E-01-.877316710E-04    3
 .551440390E-07-.141557690E-10 .392169020E+05 .371208190E+02                   4
C6H5OH                  C   6H   6O   1     G    300.00   4000.00 1000.00      1
 .141552427E+02 .199350340E-01-.718219540E-05 .116229002E-08-.697147483E-13    2
-.181287441E+05-.517984911E+02-.290978575E+00 .408562397E-01 .242829425E-04    3
-.714477617E-07 .346002146E-10-.134129780E+05 .268745637E+02                   4
C6H6O3                  C   6H   6O   3     G    300.00   4000.00 1382.00      1
 .193892545E+02 .186134462E-01-.631148097E-05 .975462374E-09-.564561412E-13    2
-.492678935E+05-.716786498E+02 .598814621E+00 .618493802E-01-.438009436E-04    3
 .155531333E-07-.220506530E-11-.427313109E+05 .293828012E+02                   4
CYC6H8                  C   6H   8          G    300.00   4000.00 1384.00      1
 .167797183E+02 .200748305E-01-.710732570E-05 .112925397E-08-.665827513E-13    2
 .222453062E+04-.729120687E+02-.719572313E+01 .780676798E-01-.620002183E-04    3
 .253310854E-07-.423684696E-11 .104082650E+05 .552451233E+02                   4
!C5H5CH3                   C   6H   8          G    300.00   4000.00 1399.00      1 !polimi
! .154352848E+02 .199801707E-01-.680270423E-05 .105349633E-08-.610336727E-13    2
! .447456576E+04-.636393642E+02-.665320026E+01 .744640477E-01-.582864186E-04    3
! .231603543E-07-.369017129E-11 .117669311E+05 .538162769E+02                   4
C5H5CH3                 C   6H   8          G    300.00   4000.00 1000.00      1 ! Burcat kik 5-Methyl-1,3-CYCLOPENTADIENE
 1.12002638E+01 2.50104924E-02-8.94914815E-06 1.44109704E-09-8.61256818E-14    2
 7.66096956E+03-3.68265351E+01 2.93206487E+00 1.12663266E-02 9.41193663E-05    3
-1.36178031E-07 5.64768524E-11 1.15372662E+04 1.42303662E+01 1.35013031E+04    4
!C5H5CH3                   C   6H   8          G    300.00   4000.00 1399.00      1 ! Burcat kik  3-METHYL-1,3-CYCLOPENTADIENE
! 1.11438571E+01 2.51265706E-02-9.00536078E-06 1.45167109E-09-8.68188102E-14    2
! 6.15685018E+03-3.61900531E+01 3.15023799E+00 1.30929547E-02 8.49819174E-05    3
!-1.23780433E-07 5.11852420E-11 9.89179835E+03 1.29939079E+01 1.19433443E+04    4
DMF                     C   6H   8O   1     G    300.00   4000.00 1000.00      1
 .117792073E+02 .285086757E-01-.111333319E-04 .199173491E-08-.133982691E-12    2
-.211130695E+05-.374257400E+02 .803526924E+00 .443305994E-01 .419434116E-05    3
-.349560898E-07 .165826978E-10-.172836857E+05 .230189579E+02                   4
C6H8O4                  C   6H   8O   4     G    300.00   4000.00 1398.00      1
 .245389912E+02 .222706283E-01-.773806446E-05 .121423501E-08-.709771757E-13    2
-.816610603E+05-.100550137E+03-.460104207E+01 .100736116E+00-.905484350E-04    3
 .413812870E-07-.752102026E-11-.725801173E+05 .522649333E+02                   4
CYC6H10                 C   6H  10          G    300.00   4000.00 1388.00      1
 .164687940E+02 .250464584E-01-.873323457E-05 .137353265E-08-.804138942E-13    2
-.977694533E+04-.696690108E+02-.607599781E+01 .751138370E-01-.506516889E-04    3
 .171683701E-07-.235089637E-11-.166592755E+04 .523699408E+02                   4
C6H10                   C   6H  10          G    300.00   4000.00 1413.00      1
 .160456030E+02 .234774145E-01-.785797929E-05 .120200542E-08-.690100029E-13    2
 .211899382E+04-.588452460E+02-.101375402E+01 .638242808E-01-.440653860E-04    3
 .158295163E-07-.230830701E-11 .794033696E+04 .325056094E+02                   4
CYC6H10-O-14            C   6H  10O   1     G    300.00   4000.00 1381.00      1
 .208569012E+02 .251723586E-01-.898344923E-05 .143508332E-08-.849382249E-13    2
-.384586302E+05-.102070819E+03-.138345764E+02 .100994913E+00-.688346635E-04    3
 .212451763E-07-.229797219E-11-.260978348E+05 .857505804E+02                   4
C5H9CHO                 C   6H  10O   1     G    300.00   4000.00 1000.00      1
 .555649280E+01 .338399710E-01-.129908190E-04 .225842790E-08-.147803790E-12    2
-.155583360E+05 .376697540E+01 .117554640E+01 .506138280E-01-.305173360E-04    3
 .629100420E-08 .920183740E-12-.149438880E+05 .244076960E+02                   4
CYC6H10-ONE             C   6H  10O   1     G    300.00   4000.00 1382.00      1
 .189587175E+02 .263606964E-01-.929344737E-05 .147257311E-08-.866645349E-13    2
-.391424596E+05-.835594309E+02-.541298687E+01 .749581025E-01-.429010347E-04    3
 .103686234E-07-.655858987E-12-.298390440E+05 .503037294E+02                   4
CYC6H10-O-12            C   6H  10O   1     G    300.00   4000.00 1388.00      1
 .211309516E+02 .245922161E-01-.870218393E-05 .138238722E-08-.815033630E-13    2
-.270082298E+05-.100017882E+03-.102441734E+02 .947119743E-01-.662992744E-04    3
 .218368996E-07-.269065692E-11-.159562249E+05 .693449458E+02                   4
CYC6H10-O-13            C   6H  10O   1     G    300.00   4000.00 1384.00      1
 .209040427E+02 .249694592E-01-.887525958E-05 .141404459E-08-.835397954E-13    2
-.281106427E+05-.100684615E+03-.120242065E+02 .974927920E-01-.669797836E-04    3
 .211938876E-07-.242310206E-11-.164176421E+05 .774198780E+02                   4
HEXENAL                 C   6H  10O   1     G    300.00   4000.00 1000.00      1
 .163810350E+02 .253163710E-01-.817955520E-05 .126084900E-08-.759870140E-13    2
-.236222230E+05-.549602890E+02 .549190040E+00 .602940540E-01-.317306290E-04    3
 .455543960E-08 .102256280E-11-.184722190E+05 .298272340E+02                   4
CYC6-OQOOH-3            C   6H  10O   3     G    300.00   4000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.696293762E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .532148412E+02                   4
ALDEST                  C   6H  10O   3     G    300.00   4000.00 1384.00      1
 .212949599E+02 .266487791E-01-.898035403E-05 .137511216E-08-.789865729E-13    2
-.762788357E+05-.785214726E+02 .521237801E+01 .613142880E-01-.373337900E-04    3
 .119679719E-07-.162337383E-11-.703135588E+05 .903341827E+01                   4
CYC6-OQOOH-2            C   6H  10O   3     G    300.00   4000.00 1416.00      1
 .160913887E+02 .291196520E-01-.940602358E-05 .140488615E-08-.793370497E-13    2
-.378857796E+05-.754185099E+02-.107476916E+02 .986835275E-01-.783513685E-04    3
 .322824282E-07-.532533650E-11-.294335398E+05 .659825481E+02                   4
CYC6-OQOOH-4            C   6H  10O   3     G    300.00   4000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.703238906E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .525203269E+02                   4
C6H10O5                 C   6H  10O   5     G    300.00   4000.00 1000.00      1
 .279850422E+02 .264166682E-01-.913640739E-05 .142923991E-08-.833656585E-13    2
-.114313686E+06-.117754445E+03-.781241700E+01 .125424511E+00-.116271866E-03    3
 .544734561E-07-.100746170E-10-.103428291E+06 .690300863E+02                   4
NC6H12                  C   6H  12          G    300.00   4000.00 1000.00      1
 .186637886E+02 .209714510E-01-.310828090E-05-.686516180E-09 .160236080E-12    2
-.135910200E+05-.708905467E+02 .196862030E+01 .476562310E-01 .660153730E-05    3
-.371481730E-07 .169224630E-10-.771187890E+04 .208592300E+02                   4
CYC6H12                 C   6H  12          G    300.00   4000.00 1373.00      1
 .190852614E+02 .283866516E-01-.999547753E-05 .158256182E-08-.930877430E-13    2
-.260770569E+05-.880292959E+02-.782903355E+01 .809375102E-01-.439655186E-04    3
 .871887784E-08-.486950162E-15-.157787533E+05 .600472718E+02                   4
DIPE                    C   6H  14O   1     G    300.00   4000.00 1000.00      1
 .961994133E+01 .527564090E-01-.244349190E-04 .491563770E-08-.360965330E-12    2
-.452985516E+05-.220408754E+02-.207944820E+01 .869029220E-01-.602649600E-04    3
 .209337360E-07-.299614610E-11-.422065600E+05 .378635810E+02                   4
TAME                    C   6H  14O   1     G    300.00   4000.00 1000.00      1
 .102413361E+02 .494717450E-01-.210657300E-04 .406005360E-08-.291140680E-12    2
-.438310029E+05-.257392482E+02-.184725690E+01 .864624650E-01-.624059780E-04    3
 .241227640E-07-.391573010E-11-.407484470E+05 .356637750E+02                   4
ETBE                    C   6H  14O   1     G    300.00   4000.00 1000.00      1
 .107600227E+02 .484809450E-01-.204693300E-04 .391707780E-08-.279248340E-12    2
-.456695052E+05-.288336460E+02-.321171820E+01 .924083860E-01-.712212230E-04    3
 .295255040E-07-.509148160E-11-.421838470E+05 .417951430E+02                   4
C6H5CHO                 C   7H   6O   1     G    200.00   6000.00 1000.00      1   !Burcat MP e Kik 20/10/17
 1.56015162E+01 2.18827888E-02-8.01082769E-06 1.30962791E-09-7.91372656E-14    2
-1.20437393E+04-5.86979950E+01 1.57674040E+00 3.02180643E-02 5.99285319E-05    3
-1.09114726E-07 4.80953568E-11-6.86186490E+03 2.06412628E+01-4.71212086E+03    4
!C6H5CHO                 C   7H   6O   1     G    300.00   4000.00 1000.00      1
! .151976148E+02 .229544430E-01-.714039470E-05 .736589790E-09 .000000000E+00    2
!-.120582935E+05-.546270656E+02-.328352400E+01 .610821620E-01-.279524170E-04    3
! .190203190E-08 .000000000E+00-.599503400E+04 .449259300E+02                   4 
!C7H8                    C   7H   8          G    300.00   4000.00 1000.00      1 ! polimi
! .988928700E+01 .312351700E-01-.110466410E-04 .129795100E-08 .000000000E+00    2
! .590756417E+03-.294263546E+02-.469518200E+01 .695108030E-01-.438445020E-04    3
! .104046480E-07 .000000000E+00 .469335500E+04 .464073200E+02                   4
C7H8  Toluene     g 1/93C  7.H  8.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.29393610E+01 2.66922277E-02-9.68422041E-06 1.57392386E-09-9.46671699E-14    2
-6.76971149E+02-4.67249759E+01 1.61200102E+00 2.11179855E-02 8.53239986E-05    3
-1.32568501E-07 5.59411406E-11 4.09654820E+03 2.02969771E+01 6.03402967E+03    4
CRESOL                  C   7H   8O   1     G    300.00   4000.00 1000.00      1
 .109411883E+02 .359221340E-01-.155859930E-04 .305336930E-08-.221926260E-12    2
-.211837368E+05-.322120090E+02-.410479790E+01 .823735850E-01-.680002460E-04    3
 .287114670E-07-.487123580E-11-.173767210E+05 .440872850E+02                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   4000.00 1000.00      1
 .988928700E+01 .312351700E-01-.110466410E-04 .129795100E-08 .000000000E+00    2
-.176276686E+05-.230348046E+02-.469518200E+01 .695108030E-01-.438445020E-04    3
 .104046480E-07 .000000000E+00-.135250700E+05 .527988700E+02                   4
C6H5OCH3                C   7H   8O   1     G    300.00   4000.00 1393.00      1
 .203938728E+02 .209088165E-01-.722522263E-05 .112997840E-08-.659097524E-13    2
-.186061425E+05-.862920505E+02-.540888697E+01 .873332441E-01-.739639658E-04    3
 .320208039E-07-.556946955E-11-.102821510E+05 .500696056E+02                   4
DIMEPTD                 C   7H  12          G    300.00   4000.00 1000.00      1
 .140192352E+02 .351774100E-01-.121769020E-04 .195853870E-08-.120886390E-12    2
-.562170122E+04-.461295916E+02 .191804150E+01 .620151830E-01-.182958650E-04    3
-.181326460E-07 .113526820E-10-.217165720E+04 .175128710E+02                   4
C7DIONE                 C   7H  12O   2     G    300.00   4000.00 1676.00      1
 .218722874E+02 .369330034E-01-.137295934E-04 .226033024E-08-.136759137E-12    2
-.450225188E+05-.973652620E+02 .236568827E+01 .679632843E-01-.230649606E-04    3
-.260553450E-08 .197085207E-11-.372372626E+05 .120380792E+02                   4
KMCYC6                  C   7H  12O   3     G    300.00   4000.00 1380.00      1
 .281047951E+02 .298656134E-01-.103750111E-04 .162883933E-08-.952775107E-13    2
-.587524861E+05-.124642473E+03-.502703972E+01 .104102110E+00-.722526077E-04    3
 .243793077E-07-.320129183E-11-.470307327E+05 .542550536E+02                   4
NC7H14                  C   7H  14          G    300.00   4000.00 1390.00      1
 .206190401E+02 .314852991E-01-.107162057E-04 .165827662E-08-.959911785E-13    2
-.196710875E+05-.822507478E+02-.116533279E+01 .790439806E-01-.496101666E-04    3
 .158569009E-07-.205346433E-11-.117362359E+05 .359871070E+02                   4
MCYC6                   C   7H  14          G    300.00   4000.00 1381.00      1
 .220211359E+02 .332076617E-01-.115857900E-04 .182324838E-08-.106797390E-12    2
-.311719553E+05-.103211614E+03-.890848850E+01 .969226774E-01-.576085500E-04    3
 .148743771E-07-.111357720E-11-.196669630E+05 .657804644E+02                   4
C7KETONE                C   7H  14O   1     G    300.00   4000.00 1385.00      1
 .232764710E+02 .323525773E-01-.112350736E-04 .176201535E-08-.102947816E-12    2
-.448556012E+05-.937710798E+02-.318897678E+00 .833005520E-01-.531219909E-04    3
 .175654519E-07-.244145064E-11-.361006378E+05 .346722541E+02                   4
NC7H14O                 C   7H  14O   1     G    300.00   4000.00 1397.00      1
 .231122557E+02 .333659362E-01-.114966228E-04 .179372703E-08-.104427245E-12    2
-.438636425E+05-.993466782E+02-.767475343E+01 .108451023E+00-.827531084E-04    3
 .330380469E-07-.541492429E-11-.334640974E+05 .649157213E+02                   4
NC7H13OOH               C   7H  14O   2     G    300.00   4000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
NC7-OQOOH               C   7H  14O   3     G    300.00   4000.00 1387.00      1
 .288332529E+02 .320168096E-01-.111508456E-04 .175226159E-08-.102520451E-12    2
-.622309509E+05-.116187714E+03 .152936692E+01 .958173466E-01-.696688520E-04    3
 .269540382E-07-.438728126E-11-.526003608E+05 .306986714E+02                   4
NC7H16                  C   7H  16          G    300.00   4000.00 1000.00      1
 .205103125E+02 .346389640E-01-.107743740E-04 .160399760E-08-.937017530E-13    2
-.326499224E+05-.807081180E+02-.679531340E+00 .810756760E-01-.423279310E-04    3
 .697965770E-08 .837326950E-12-.256907030E+05 .329815600E+02                   4
NC7H15OOH               C   7H  16O   2     G    300.00   4000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
C8H2                    C   8H   2          G    300.00   4000.00 1000.00      1
 .156802100E+02 .111546100E-01-.372437300E-05 .519789100E-09-.237555000E-13    2
 .108112300E+06-.557143700E+02 .463042700E+01 .393708000E-01-.114803500E-04    3
-.256221400E-07 .167079100E-10 .110828500E+06 .807742500E+00                   4
!C6H5C2H                 C   8H   6          G    300.00   4000.00 1399.00      1 !Polimi
! .190886756E+02 .170819066E-01-.559393248E-05 .845345947E-09-.482537486E-13    2
! .280711996E+05-.790035627E+02-.377007730E+01 .792380003E-01-.711832819E-04    3
! .324077613E-07-.583009863E-11 .350595597E+05 .405332699E+02                   4
C6H5C2H  C6H5CCH  T12/06C  8.H  6.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.63582907E+01 2.11974105E-02-7.65817215E-06 1.24134505E-09-7.45327960E-14    2
 3.10375340E+04-6.22520227E+01-2.74707918E+00 7.78284438E-02-6.69709932E-05    3
 2.37972496E-08-8.43279765E-13 3.61131008E+04 3.54221257E+01 3.82082350E+04    4
BZFUR                   C   8H   6O   1     G    300.00   4000.00 1000.00      1
 .161267559E+02 .242942790E-01-.882919089E-05 .143722155E-08-.865592465E-13    2
-.574867958E+04-.640564836E+02-.785221476E+00 .396432449E-01 .569751746E-04    3
-.114831806E-06 .519411145E-10 .215748538E+03 .302655928E+02                   4
!C6H5C2H3                C   8H   8          G    300.00   4000.00 1000.00      1 !Polimi
! .132118086E+02 .297097690E-01-.100379980E-04 .113030440E-08 .000000000E+00    2
! .112255113E+05-.452965784E+02-.314842000E+01 .733550410E-01-.482478610E-04    3
! .120551240E-07 .000000000E+00 .157685200E+05 .395339300E+02                   4
C6H5C2H3 Styrene  T12/10C  8.H  8.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.55820120E+01 2.66093018E-02-9.56144870E-06 1.54378205E-09-9.24814823E-14    2
 1.03197319E+04-5.98622481E+01 1.12656107E+00 3.17044880E-02 7.38511452E-05    3
-1.29131757E-07 5.65307288E-11 1.57676346E+04 2.25936971E+01 1.79366548E+04    4
!C6H5C2H5                C   8H  10          G    300.00   4000.00 1000.00      1 !Polimi
! .123967254E+02 .365194120E-01-.128125900E-04 .149467160E-08 .000000000E+00    2
!-.304290347E+04-.409211516E+02-.458801200E+01 .813929890E-01-.516055260E-04    3
! .123987680E-07 .000000000E+00 .171000000E+04 .472934500E+02                   4
C6H5C2H5          A11/04C  8.H 10.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.56901336E+01 3.23663075E-02-1.16864578E-05 1.88989562E-09-1.13201791E-13    2
-4.38669907E+03-6.04442403E+01 1.24076722E+00 3.59132829E-02 7.54222474E-05    3
-1.31904301E-07 5.74746803E-11 1.18391719E+03 2.24682133E+01 3.58290266E+03    4
!XYLENE                  C   8H  10          G    300.00   4000.00 1000.00      1 ! polimi
! .104572604E+02 .403200160E-01-.145441770E-04 .173870560E-08 .000000000E+00    2
!-.392485555E+04-.316838798E+02-.365621300E+01 .742185790E-01-.400008720E-04    3
! .741031100E-08 .000000000E+00 .307000000E+03 .427477900E+02                   4
XYLENE  o-Di-Met  T 9/13C  8.H 10.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.38533968E+01 3.30836404E-02-1.18974456E-05 1.92231652E-09-1.15153932E-13    2
-5.17475507E+03-5.00163449E+01 2.96890501E+00 2.10981093E-02 9.87221885E-05    3
-1.46214604E-07 6.02721557E-11-2.13940788E+02 1.61289213E+01 2.22069515E+03    4
C8H10O3                 C   8H  10O   3     G    300.00   4000.00 1280.00      1
 .386588321E+02 .317536134E-02 .740594019E-05-.343506103E-08 .445199316E-12    2
-.597114304E+05-.165594980E+03 .580160876E+00 .872417598E-01-.555691469E-04    3
 .111625328E-07 .157789482E-11-.515704990E+05 .289562016E+02                   4
UME7                    C   8H  14O   2     G    300.00   4000.00 1386.00      1
 .274195251E+02 .331653074E-01-.112369879E-04 .173174767E-08-.999867016E-13    2
-.597230517E+05-.112624254E+03 .202528941E+01 .898844344E-01-.593620598E-04    3
 .203016355E-07-.286718129E-11-.505953610E+05 .247655861E+02                   4
IC8H16                  C   8H  16          G    300.00   4000.00 1000.00      1
 .159403331E+02 .467083530E-01-.162445520E-04 .262105430E-08-.162114790E-12    2
-.212288474E+05-.575000710E+02-.188446240E+01 .875446570E-01-.337527930E-04    3
-.140196880E-07 .109753600E-10-.160534330E+05 .363096160E+02                   4
IC8H16O                 C   8H  16O   1     G    300.00   4000.00 1400.00      1
 .286870453E+02 .350973257E-01-.120318626E-04 .187165307E-08-.108763411E-12    2
-.489758985E+05-.130519447E+03-.811336944E+01 .120858100E+00-.869108786E-04    3
 .308943900E-07-.431018679E-11-.363657206E+05 .668763983E+02                   4
IC8-OQOOH               C   8H  16O   3     G    300.00   4000.00 1395.00      1
 .329665839E+02 .352889373E-01-.121856584E-04 .190423031E-08-.110989507E-12    2
-.686224367E+05-.138776314E+03 .233137835E+00 .110643301E+00-.779138892E-04    3
 .277663606E-07-.398875833E-11-.571903320E+05 .373387625E+02                   4
IC8H18                  C   8H  18          G    300.00   4000.00 1000.00      1
 .175409498E+02 .499242880E-01-.172020170E-04 .275518900E-08-.169419330E-12    2
-.363533756E+05-.670046390E+02-.203218650E+01 .946845260E-01-.357433050E-04    3
-.165946760E-07 .125346320E-10-.306832730E+05 .359861450E+02                   4
!INDENE                  C   9H   8          G    300.00   4000.00 1000.00      1 !polimi
! .129942100E+02 .345035980E-01-.119473340E-04 .137705200E-08 .000000000E+00    2
! .128398488E+05-.468095535E+02-.565650900E+01 .835992990E-01-.541865810E-04    3
! .131713170E-07 .000000000E+00 .180739000E+05 .501175500E+02                   4
INDENE            T 9/96C  9.H  8.   0.   0.G   200.000  6000.000  1000.       1 !Burcat kik
 1.73186757E+01 2.89827586E-02-1.06050551E-05 1.73345448E-09-1.04679146E-13    2
 1.11514275E+04-7.15553836E+01-6.81899560E-01 4.16587045E-02 7.07413209E-05    3
-1.34308856E-07 5.99158843E-11 1.77050360E+04 2.97813474E+01 1.97411898E+04    4
C9H10O2                 C   9H  10O   2     G    300.00   4000.00 1400.00      1
 .279893805E+02 .257305292E-01-.858901356E-05 .131357222E-08-.754726372E-13    2
-.378460988E+05-.119703580E+03-.219761532E+01 .995964750E-01-.769418656E-04    3
 .296736479E-07-.451992280E-11-.279092089E+05 .408797910E+02                   4
TMBENZ                  C   9H  12          G    300.00   4000.00 1383.00      1
 .215885246E+02 .321229102E-01-.110727239E-04 .172825742E-08-.100649304E-12    2
-.136169019E+05-.914142733E+02-.173308850E+01 .786049041E-01-.431048197E-04    3
 .100745302E-07-.585489308E-12-.471446607E+04 .366811038E+02                   4
NPBENZ                  C   9H  12          G    300.00   4000.00 1395.00      1
 .234758956E+02 .300348225E-01-.102493106E-04 .158931255E-08-.921475616E-13    2
-.109980792E+05-.102092892E+03-.597461242E+01 .101439137E+00-.768408376E-04    3
 .299742828E-07-.474668103E-11-.108882285E+04 .550543799E+02                   4
C7H15COCHO              C   9H  16O   2     G    300.00   4000.00 1387.00      1
 .303225194E+02 .381334789E-01-.128450948E-04 .197085647E-08-.113456990E-12    2
-.668175594E+05-.126355483E+03-.229351926E+00 .108754598E+00-.755330139E-04    3
 .275093508E-07-.415197146E-11-.560981532E+05 .380532571E+02                   4
ALD9                    C   9H  18O   1     G    300.00   4000.00 1000.00      1
 .106561750E+02 .676363860E-01-.253129890E-04 .432392120E-08-.279580530E-12    2
-.437018400E+05-.154058910E+02-.276341620E+00 .105894390E+00-.646322300E-04    3
 .149734250E-07 .101003800E-11-.417122110E+05 .376426280E+02                   4
C10H8                   C  10H   8          G    300.00   4000.00 1401.00      1
 .234023214E+02 .242434427E-01-.836282016E-05 .130620111E-08-.761153748E-13    2
 .651941329E+04-.107433208E+03-.883645988E+01 .109300567E+00-.955200914E-04    3
 .421647669E-07-.739851710E-11 .166533366E+05 .621064766E+02                   4
C10H7OH                 C  10H   8O   1     G    300.00   4000.00 1394.00      1
 .262017858E+02 .245473904E-01-.859268465E-05 .135522543E-08-.795056830E-13    2
-.158010339E+05-.119344614E+03-.322687986E+01 .931430619E-01-.687932451E-04    3
 .249753868E-07-.357353464E-11-.568766282E+04 .385570421E+02                   4
C9H9              -----0H   9C   9          G     300.0    5000.0  1000.0    0 1  !AN 2100 from Jin et al 2019; to be rescaled wrt steady state branching of C9H9-1,C9H9-2,A1C3H4
   1.58195435E1  3.45357901E-2 -1.36013494E-5   2.4480452E-9-1.65409696E-13    2
   1.62783704E4  -6.19015515E1   -7.0786938E0  9.13681374E-2 -5.31256325E-5    3
-8.66380926E-10 8.66347995E-12   2.29720325E4   5.80700378E1                   4
FC10H10                 H  10C  10          G   290.000  2500.000  997.76      1  !AN 2100 from Long et al 2018; ONLY ISOMER T1A. IRRELEVANT BECAUSE NO EQ. REACTIONS INCLUDED
 3.74069224E+00 7.54937065E-02-4.97910050E-05 1.64156284E-08-2.14692831E-12    2
 3.06016191E+04 1.60008660E+00-4.08179268E+00 8.55612763E-02-3.29153684E-05    3
-1.62487375E-08 1.13967163E-11 3.32224694E+04 4.46327208E+01                   4
FC10H10O                H  10C  10O   1     G   290.000  2500.000  997.76      1  ! LPM SAME AS C10H10, WRONG BUT TEMPORARY
 3.74069224E+00 7.54937065E-02-4.97910050E-05 1.64156284E-08-2.14692831E-12    2
 3.06016191E+04 1.60008660E+00-4.08179268E+00 8.55612763E-02-3.29153684E-05    3
-1.62487375E-08 1.13967163E-11 3.32224694E+04 4.46327208E+01                   4
!C10H10                  C  10H  10          G    300.00   4000.00 2043.00      1
! .196465049E+02 .362867673E-01-.135117921E-04 .222712581E-08-.134868100E-12    2
! .466515480E+04-.883925826E+02-.975555457E+01 .989343734E-01-.593843991E-04    3
! .154882804E-07-.129445409E-11 .148791325E+05 .708155586E+02                   4
C10H10                  C  10H  10          G    200.00   6000.00 1000.00      1  !AN 2100 from Long et al 2018 - most stable isomer from lumping
 1.92211178E+01 3.51247274E-02-1.27719042E-05 2.07903232E-09-1.25191968E-13    2
 4.39595221E+03-8.19390283E+01-1.92135165E-01 4.50394780E-02 8.64482370E-05    3
-1.56640588E-07 6.88727900E-11 1.16587583E+04 2.82951960E+01 1.40900666E+04    4
TETRALIN                C  10H  12          G    300.00   4000.00 1393.00      1
 .259510150E+02 .311178636E-01-.105072610E-04 .161945272E-08-.935513420E-13    2
-.106963510E+05-.121999608E+03-.103201470E+02 .118533935E+00-.903074920E-04    3
 .343768814E-07-.519161790E-11 .142964373E+04 .715127353E+02                   4
DCYC5                   C  10H  16          G    300.00   4000.00 1396.00      1
 .273482865E+02 .461538793E-01-.158755646E-04 .247442795E-08-.143965250E-12    2
-.380245063E+05-.136978542E+03-.149885463E+02 .144180968E+00-.101905712E-03    3
 .365256640E-07-.527588038E-11-.233132452E+05 .905738933E+02                   4
KHDECA                  C  10H  16O   3     G    300.00   4000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.703238906E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .525203269E+02                   4
DECALIN                 C  10H  18          G    300.00   4000.00 1396.00      1
 .273482865E+02 .461538793E-01-.158755646E-04 .247442795E-08-.143965250E-12    2
-.380245063E+05-.136978542E+03-.149885463E+02 .144180968E+00-.101905712E-03    3
 .365256640E-07-.527588038E-11-.233132452E+05 .905738933E+02                   4
ODECAL                  C  10H  18          G    300.00   4000.00 1383.00      1
 .304308606E+02 .423969327E-01-.145305017E-04 .226051483E-08-.131385276E-12    2
-.274622725E+05-.143201137E+03-.921337866E+01 .127293330E+00-.797537373E-04    3
 .229874961E-07-.227548927E-11-.131010829E+05 .721555536E+02                   4
MEALD9                  C  10H  18O   3     G    300.00   4000.00 1000.00      1
-.690383480E+01 .109133900E+00-.458269710E-04 .848431460E-08-.580474200E-12    2
-.758799840E+05 .927347110E+02-.868940000E+00 .130857110E+00-.927276920E-04    3
 .252031600E-07 .168027310E-11-.817747730E+05 .466361500E+02                   4
NC10H20                 C  10H  20          G    300.00   4000.00 1390.00      1
 .306417045E+02 .444757412E-01-.152579717E-04 .237363570E-08-.137907421E-12    2
-.321647483E+05-.129750528E+03-.253770965E+01 .118319727E+00-.776112696E-04    3
 .262647573E-07-.366153318E-11-.202029921E+05 .498650630E+02                   4
NC10MOOH                C  10H  20O   2     G    300.00   4000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
NC10-OQOOH              C  10H  20O   3     G    300.00   4000.00 1390.00      1
 .373427699E+02 .457774433E-01-.156578702E-04 .243101177E-08-.141046271E-12    2
-.740262240E+05-.156527917E+03 .209018845E+01 .128739739E+00-.918467610E-04    3
 .350282382E-07-.560696315E-11-.617151278E+05 .328016208E+02                   4
NC10H22                 C  10H  22          G    300.00   4000.00 1391.00      1
 .319882239E+02 .477244922E-01-.162276391E-04 .250963259E-08-.145215772E-12    2
-.466392840E+05-.137615344E+03-.208416969E+01 .122535012E+00-.776815739E-04    3
 .249834877E-07-.323548038E-11-.343021863E+05 .471147911E+02                   4
!C10H7CHO                C  11H   8O   1     G    300.00   4000.00 1391.00      1 !Polimi
! .276532029E+02 .258287942E-01-.902879433E-05 .142281038E-08-.834251834E-13    2
!-.106453206E+05-.124981465E+03-.108527081E+01 .881681978E-01-.575973932E-04    3
! .170999043E-07-.173813923E-11-.356369995E+03 .307785222E+02                   4
C10H7CHO          T 7/98C  11H   8O   1    0G   200.000  6000.000 1000.        1 !Burcat kik
 2.42593357E+01 3.16036997E-02-1.18467358E-05 1.96728679E-09-1.20096869E-13    2
-7.83388781E+03-1.07718994E+02-3.75140208E-01 6.11007395E-02 4.92528177E-05    3
-1.17296000E-07 5.31810720E-11 8.41138142E+02 2.88322573E+01 3.67348166E+03    4
!C10H7CH3                C  11H  10          G    300.00   4000.00 1394.00      1 !Polimi
! .269623579E+02 .288172394E-01-.100254209E-04 .157466721E-08-.921126923E-13    2
! .586670370E+03-.125206708E+03-.798962224E+01 .117448428E+00-.976360478E-04    3
! .414932114E-07-.710609396E-11 .120022223E+05 .599922187E+02                   4
C10H7CH3          T 7/98C  11H  10    0    0G   200.000  6000.000 1000.        1 !Burcat kik
 2.17939213E+01 3.60214098E-02-1.33228698E-05 2.19304403E-09-1.33071380E-13    2
 3.16261439E+03-9.48675403E+01-1.03043715E+00 6.03358177E-02 5.45655719E-05    3
-1.22769251E-07 5.54507327E-11 1.13241014E+04 3.22970611E+01 1.39642625E+04    4
CH3C10H6OH              C  11H  10O   1     G    300.00   4000.00 1392.00      1
 .281549167E+02 .299236572E-01-.104056239E-04 .163381420E-08-.955470229E-13    2
-.208064399E+05-.126965793E+03-.171335238E+01 .970093442E-01-.665430499E-04    3
 .223717851E-07-.293871610E-11-.102462828E+05 .342637221E+02                   4
C11H12O4                C  11H  12O   4     G    300.00   4000.00 1398.00      1
 .495886732E+02 .844753396E-02 .385179844E-05-.232491508E-08 .315199759E-12    2
-.164047630E+05-.193448260E+03 .542487420E+01 .999122905E-01-.513976516E-04    3
-.430175388E-08 .876106788E-11-.572347637E+04 .356171545E+02                   4
UME10                   C  11H  20O   2     G    300.00   4000.00 1384.00      1
 .374112533E+02 .458948435E-01-.156057696E-04 .241315080E-08-.139673864E-12    2
-.736971925E+05-.162545741E+03 .937241013E+00 .126885097E+00-.836053178E-04    3
 .282312118E-07-.390359926E-11-.605539595E+05 .349335674E+02                   4
ETEROMD                 C  11H  20O   3     G    300.00   4000.00 1386.00      1
 .418053606E+02 .443798286E-01-.151698489E-04 .235874245E-08-.137104681E-12    2
-.896960798E+05-.186388223E+03-.869108022E+00 .143689897E+00-.103700029E-03    3
 .384483018E-07-.582555005E-11-.748416098E+05 .429341731E+02                   4
MDKETO                  C  11H  20O   5     G    300.00   4000.00 1391.00      1
 .435827467E+02 .471875465E-01-.155121189E-04 .235632808E-08-.134947249E-12    2
-.114156459E+06-.184940808E+03 .336575533E+01 .147442203E+00-.113482823E-03    3
 .468018272E-07-.796034235E-11-.100759720E+06 .289177372E+02                   4
MD                      C  11H  22O   2     G    300.00   4000.00 1382.00      1
 .393230373E+02 .488368389E-01-.166923510E-04 .259065840E-08-.150309877E-12    2
-.885441006E+05-.173932688E+03 .176901386E+01 .129360919E+00-.808243357E-04    3
 .251676921E-07-.312062272E-11-.747104475E+05 .304352079E+02                   4
!C12H8                   C  12H   8          G    300.00   4000.00 1000.00      1 !polimi
! .213682716E+02 .324830670E-01-.101214580E-04 .104613640E-08 .000000000E+00    2
! .210494631E+05-.924787980E+02-.672892800E+01 .106967800E+00-.747993040E-04    3
! .193364490E-07 .000000000E+00 .288910000E+05 .533672000E+02                   4
C12H8 Acenaphtyl  T01/08C 12.H  8.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 2.15561639E+01 3.31444907E-02-1.20903392E-05 1.97278991E-09-1.19007513E-13    2
 2.07186570E+04-9.76752478E+01-2.14921587E+00 5.89101361E-02 6.42492047E-05    3
-1.41293714E-07 6.47476866E-11 2.89379865E+04 3.36791245E+01 3.12345526E+04    4
DIBZFUR                 C  12H   8O   1     G    300.00   4000.00 1000.00      1
 .238928699E+02 .342239370E-01-.125916314E-04 .206592304E-08-.125089220E-12    2
-.481449779E+04-.107327684E+03-.194754604E+01 .663215475E-01 .555418713E-04    3
-.135401425E-06 .629515620E-10 .401745217E+04 .350605098E+02                   4
!BIPHENYL                C  12H  10          G    300.00   4000.00 1000.00      1 !polimi
! .214890352E+02 .375797860E-01-.121080230E-04 .129882780E-08 .000000000E+00    2
! .115420788E+05-.916763235E+02-.783196500E+01 .114327200E+00-.776398370E-04    3
! .194042280E-07 .000000000E+00 .198069600E+05 .608493300E+02                   4
BIPHENYL          g 8/00C 12.H 10.   0.   0.G   200.000  6000.000 1000.00      1 !Burcat kik
 2.28963620E+01 3.68453189E-02-1.35016357E-05 2.20802787E-09-1.33358137E-13    2
 1.07395923E+04-1.00509573E+02 1.94600056E-01 5.35259888E-02 8.55000841E-05    3
-1.63903525E-07 7.29975666E-11 1.90021492E+04 2.72148992E+01 2.19050792E+04    4
C6H5OC6H5               C  12H  10O   1     G    300.00   4000.00 1000.00      1
 .283319364E+02 .317670352E-01-.107447484E-04 .165690065E-08-.957158914E-13    2
-.789446240E+04-.127230446E+03-.865410063E+01 .124988347E+00-.100933530E-03    3
 .413234204E-07-.675938299E-11 .409381103E+04 .686981333E+02                   4
C12H18                  C  12H  18          G    300.00   4000.00 1000.00      1
 .938665800E+02 .198595000E-01-.295692400E-05 .245328200E-09-.917006600E-14    2
-.897187500E+05-.457207000E+03 .374918500E+01 .185852000E+00-.868236800E-04    3
 .615957800E-08 .205893500E-11-.565341800E+05 .387544400E+02                   4
C12H22                  C  12H  22          G    300.00   4000.00 1392.00      1
 .362943970E+02 .488870789E-01-.165740715E-04 .255852468E-08-.147868438E-12    2
-.229987583E+05-.159907963E+03-.329755440E+01 .140713318E+00-.978288195E-04    3
 .352594898E-07-.520523450E-11-.920475977E+04 .529246931E+02                   4
NC12-OQOOH              C  12H  24O   3     G    300.00   4000.00 1678.00      1
 .447068212E+02 .522272795E-01-.195350799E-04 .322923457E-08-.195935332E-12    2
-.818914807E+05-.192299360E+03 .877388676E+01 .119113497E+00-.561329021E-04    3
 .677643630E-08 .106366869E-11-.685051188E+05 .572134782E+01                   4
NC12H26                 C  12H  26          G    300.00   4000.00 1391.00      1
 .385099212E+02 .563550048E-01-.191493200E-04 .296024862E-08-.171244150E-12    2
-.548849270E+05-.169785166E+03-.262181594E+01 .147237711E+00-.943970271E-04    3
 .307441268E-07-.403602230E-11-.400654253E+05 .529882396E+02                   4
!FLUORENE                C  13H  10          G    300.00   4000.00 1000.00      1 !Polimi
! .231612871E+02 .392128530E-01-.125431510E-04 .133503890E-08 .000000000E+00    2
! .123102892E+05-.103717257E+03-.112092800E+02 .129847800E+00-.907013380E-04    3
! .232288460E-07 .000000000E+00 .219426600E+05 .748524200E+02                   4
FLUORENE          T11/07C 13.H 10.   0.   0.G   200.000  6000.000  1000.00     1 !Burcat kik
 2.33961594E+01 3.76272122E-02-1.37117389E-05 2.24351896E-09-1.35502173E-13    2
 9.60546553E+03-1.04754427E+02-1.08010254E+00 5.81364450E-02 8.71414836E-05    3
-1.72419903E-07 7.76417263E-11 1.83197800E+04 3.21625902E+01 2.10475422E+04    4
!C6H5CH2C6H5             C  13H  12          G    300.00   4000.00 1000.00      1 !polimi
! .185418955E+02 .513343070E-01-.178726910E-04 .207043850E-08 .000000000E+00    2
! .668552054E+04-.690121392E+02-.940899900E+01 .125451300E+00-.822539730E-04    3
! .202856220E-07 .000000000E+00 .144845500E+05 .760677200E+02                   4
C6H5CH2C6H5       T10/13C 13.H 12.   0.   0.G   200.000  6000.000  1000.0      1 !Burcat kik MeBiPhenyl
 2.33823671E+01 4.36035134E-02-1.59318261E-05 2.59973976E-09-1.56760199E-13    2
 7.84267591E+03-1.00997944E+02 1.70749233E+00 3.70722686E-02 1.53928694E-04    3
-2.41954650E-07 1.02743229E-10 1.67215993E+04 2.61209040E+01 1.98087440E+04    4
ALDINS                  C  13H  20O   1     G    300.00   4000.00 1000.00      1
 .938665800E+02 .198595000E-01-.295692400E-05 .245328200E-09-.917006600E-14    2
-.897187500E+05-.457207000E+03 .374918500E+01 .185852000E+00-.868236800E-04    3
 .615957800E-08 .205893500E-11-.565341800E+05 .387544400E+02                   4
U2ME12                  C  13H  22O   2     G    300.00   4000.00 1391.00      1
 .422353117E+02 .524987045E-01-.181261023E-04 .283174793E-08-.165001495E-12    2
-.676968189E+05-.186270028E+03 .679798314E-01 .152530074E+00-.111376081E-03    3
 .435663556E-07-.715842617E-11-.529996239E+05 .399987338E+02                   4
MEALDU12                C  13H  22O   3     G    300.00   4000.00 1000.00      1
 .102076680E+02 .102462700E+00-.400200840E-04 .704170850E-08-.464730410E-12    2
-.764049450E+05 .447871400E+01-.148239800E+01 .157342330E+00-.103758050E-03    3
 .246418600E-07 .237571010E-11-.758768280E+05 .556433530E+02                   4
!C14H10                  C  14H  10          G    300.00   4000.00 1000.00      1 !polimi
! .255171870E+02 .393727940E-01-.123155080E-04 .127852800E-08 .000000000E+00    2
! .131224037E+05-.115618425E+03-.909474100E+01 .131333800E+00-.924017290E-04    3
! .240156710E-07 .000000000E+00 .227649500E+05 .639753600E+02                   4
C14H10  Phenanth  T 6/12C 14.H 10.   0.   0.G   200.000  6000.000  1000.00     1 ! Burcat kik
 2.66042825E+01 3.97675990E-02-1.45710303E-05 2.38414417E-09-1.44083321E-13    2
 1.15427370E+04-1.22473909E+02-3.36413181E+00 8.50677802E-02 3.75500017E-05    3
-1.26667049E-07 6.14543114E-11 2.14305029E+04 4.07973319E+01 2.43189316E+04    4
!C6H5C2H4C6H5            C  14H  14          G    300.00   4000.00 1000.00      1 !polimi
! .183724857E+02 .606470630E-01-.215506390E-04 .254284330E-08 .000000000E+00    2
! .518516081E+04-.659251182E+02-.814781700E+01 .130620600E+00-.819367560E-04    3
! .194757260E-07 .000000000E+00 .126141800E+05 .718458700E+02                   4
!C6H5C2H4C6H5      T 5/04C 14.H 14.   0.   0.G   200.000  6000.000  1000.00     1 !Burcat kik
! 2.65979897E+01 4.68689340E-02-1.69056103E-05 2.73737090E-09-1.64235887E-13    2
! 3.18810786E+03-1.14827874E+02 1.30521842E+00 5.76220698E-02 1.22418244E-04    3
!-2.18120750E-07 9.59096665E-11 1.26627763E+04 2.90742354E+01 1.63088384E+04    4
C6H5C2H4C6H5            C  14H  14O   0    0G   300.00   3000.00  1000.00      1 
 0.72920350E+01 0.92502000E-01-0.51686410E-04 0.13627090E-07-0.13811480E-11    2                      
 0.10316730E+05-0.11327380E+02-0.13889580E+02 0.17209840E+00-0.17006600E-03    3                      
 0.96018880E-07-0.23732530E-10 0.15032340E+05 0.92707360E+02                   4
!C16H10                  C  16H  10          G    300.00   4000.00 1000.00      1 !polimi
! .290747022E+02 .412337670E-01-.126077060E-04 .127453580E-08 .000000000E+00    2
! .141687238E+05-.136431347E+03-.106811200E+02 .146535400E+00-.103943520E-03    3
! .270645390E-07 .000000000E+00 .252715000E+05 .699617500E+02                   4
C16H10 Pyrene     T 6/12C 16.H 10.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 2.99100370E+01 4.26680281E-02-1.57338134E-05 2.58516829E-09-1.56679506E-13    2
 1.27624176E+04-1.41870304E+02-4.04244612E+00 9.15520165E-02 5.14380972E-05    3
-1.52760613E-07 7.30856860E-11 2.40702419E+04 4.36665325E+01 2.71212615E+04    4
C18H10                  C  18H  10          G    300.00   3500.00 1430.00      1 !test C18H10=C16H10+(C16H10-C14H10)
 3.55205969e+01 2.97059226e-02-5.18577408e-06-7.74976601e-10 2.05764301e-13    2
 1.13998034e+04-1.72584653e+02-1.43149515e+01 1.69106058e-01-1.51409692e-04    3
 6.73946823e-08-1.17120082e-11 2.56527702e+04 8.56679628e+01                   4
!C18H10                  C 18.H 10.          G    300.00  4000.00  1000.00      1 !  KS 1800
! 3.26322170E+01 4.3094740E-02 -1.2899904E-05  1.2705436E-09  0.0000000E+00     2
! 1.52150440E+04-1.5724427E+02 -1.2267499E+01  1.6173700E-01 -1.1548531E-04     3
! 3.01134070E-08 0.0000000E+00  2.7778050E+04  7.5948140E+01                    4
NC16-OQOOH              C  16H  32O   3     G    300.00   4000.00 1854.00      1
 .488264318E+02 .825357366E-01-.292747409E-04 .467245514E-08-.276718037E-12    2
-.942845289E+05-.205583924E+03 .138386904E+01 .198379105E+00-.134722947E-03    3
 .475955890E-07-.691333208E-11-.791319641E+05 .463051187E+02                   4
IC16-OQOOH              C  16H  32O   3     G    300.00   4000.00 1397.00      1
 .620188250E+02 .682375774E-01-.235322180E-04 .367416933E-08-.214025539E-12    2
-.107194396E+06-.296402060E+03-.700111687E+01 .236135134E+00-.181200158E-03    3
 .715715364E-07-.114883341E-10-.839739066E+05 .717765001E+02                   4
NC16H34                 C  16H  34          G    300.00   4000.00 1391.00      1
 .515593854E+02 .736064257E-01-.249888737E-04 .386085377E-08-.223263662E-12    2
-.713781425E+05-.234158439E+03-.369111950E+01 .196612966E+00-.127777824E-03    3
 .422323349E-07-.562967041E-11-.515927302E+05 .647080513E+02                   4
IC16H34                 C  16H  34          G    300.00   4000.00 1400.00      1
 .565856523E+02 .692869560E-01-.234931111E-04 .362720220E-08-.209665225E-12    2
-.820366778E+05-.276851694E+03-.107545408E+02 .233995831E+00-.178076331E-03    3
 .696956034E-07-.110282035E-10-.595981394E+05 .818346760E+02                   4
UME16                   C  17H  32O   2     G    300.00   4000.00 1000.00      1
 .333606142E+02 .106719124E+00-.429500189E-04 .790457654E-08-.546125152E-12    2
-.868236054E+05-.126816968E+03 .114310960E+02 .102101194E+00 .102480878E-03    3
-.181385357E-06 .698603588E-10-.778209017E+05 .206428096E+01                   4
ETEROMPA                C  17H  32O   3     G    300.00   4000.00 1000.00      1
 .406345250E+02 .963702350E-01-.332815250E-04 .536978820E-08-.333546480E-12    2
-.105022900E+06-.161181400E+03-.374618910E+01 .216936450E+00-.134184780E-03    3
 .217036750E-07 .800116570E-11-.930412810E+05 .677468110E+02                   4
MPA                     C  17H  34O   2     G    300.00   4000.00 1000.00      1
 .355305296E+02 .109746228E+00-.440981772E-04 .810571172E-08-.559469785E-12    2
-.102923616E+06-.145292419E+03 .117629996E+02 .108027697E+00 .103662595E-03    3
-.187190120E-06 .724616510E-10-.933306777E+05-.643066315E+01                   4
KHMLIN1                 C  19H  30O   5     G    300.00   4000.00 1843.00      1
 .597680898E+02 .832144998E-01-.302817533E-04 .491632066E-08-.294624551E-12    2
-.961002787E+05-.258440317E+03-.347354324E+01 .238348931E+00-.171810701E-03    3
 .624560833E-07-.914836595E-11-.760003616E+05 .770024622E+02                   4
MLIN1                   C  19H  32O   2     G    300.00   4000.00 1834.00      1
 .520202170E+02 .871284776E-01-.313984409E-04 .506450961E-08-.302130761E-12    2
-.727531890E+05-.226713941E+03-.298592567E+01 .218746556E+00-.148096154E-03    3
 .511216154E-07-.719451974E-11-.549290521E+05 .662774857E+02                   4
MLINO                   C  19H  34O   2     G    300.00   4000.00 1833.00      1
 .524257963E+02 .910351615E-01-.326514183E-04 .524998946E-08-.312507814E-12    2
-.869039436E+05-.227879204E+03-.158761924E+01 .219526542E+00-.145761172E-03    3
 .495347572E-07-.688636525E-11-.693288124E+05 .600962817E+02                   4
MLIN1OOH                C  19H  34O   4     G    300.00   4000.00 1833.00      1
 .524257963E+02 .910351615E-01-.326514183E-04 .524998946E-08-.312507814E-12    2
-.869039436E+05-.227879204E+03-.158761924E+01 .219526542E+00-.145761172E-03    3
 .495347572E-07-.688636525E-11-.693288124E+05 .600962817E+02                   4
MEOLE                   C  19H  36O   2     G    300.00   4000.00 1831.00      1
 .528856562E+02 .948572658E-01-.338668063E-04 .542873444E-08-.322458135E-12    2
-.101075125E+06-.229348639E+03-.267573662E+00 .220639742E+00-.143861659E-03    3
 .481699649E-07-.661786902E-11-.837166223E+05 .542791001E+02                   4
MLINOOH                 C  19H  36O   4     G    300.00   4000.00 1833.00      1
 .524257963E+02 .910351615E-01-.326514183E-04 .524998946E-08-.312507814E-12    2
-.869039436E+05-.227879204E+03-.158761924E+01 .219526542E+00-.145761172E-03    3
 .495347572E-07-.688636525E-11-.693288124E+05 .600962817E+02                   4
MSTEAKETO               C  19H  36O   5     G    300.00   4000.00 1857.00      1
 .628573476E+02 .927885184E-01-.331648431E-04 .532086973E-08-.316267196E-12    2
-.142644021E+06-.277684268E+03-.711176329E+00 .251338095E+00-.180571731E-03    3
 .664483461E-07-.990089173E-11-.122716422E+06 .585265768E+02                   4
MSTEA                   C  19H  38O   2     G    300.00   4000.00 1000.00      1
 .418174710E+02 .117959830E+00-.465265590E-04 .845319460E-08-.579171090E-12    2
-.110862900E+06-.175601040E+03 .114771030E+02 .131225240E+00 .898738730E-04    3
-.183685190E-06 .722337400E-10-.991500330E+05-.163992920E+01                   4
C24H28O4                C  24H  28O   4     G    300.00   3500.00 1080.00      1   !refitted MP
 1.29252077e+01 8.11297231e-02-4.64957369e-05 1.23575606e-08-1.22239430e-12    2
-7.66058387e+03-2.94388613e+00 3.08710528e+00 1.17567139e-01-9.71032594e-05    3
 4.35967720e-08-8.45369325e-12-5.53555376e+03 4.52764215e+01                   4
 !C24H28O4                C  24H  28O   4     G    300.00   4000.00 1398.00      1	!discontinuity highlighted
! .495886732E+02 .844753396E-02 .385179844E-05-.232491508E-08 .315199759E-12    2
!-.164047630E+05-.193448260E+03 .542487420E+01 .999122905E-01-.513976516E-04    3
!-.430175388E-08 .876106788E-11-.572347637E+04 .356171545E+02                   4
!O                       O   1               G    300.00   4000.00  700.00      1
! .854006043E+00-.488003453E-02 .104572169E-04-.522729913E-08 .771608734E-12    2
! .306893420E+05 .173763860E+02 .000000000E+00 .000000000E+00 .000000000E+00    3
! .473195502E-08-.278526775E-11 .308089029E+05 .211918689E+02                   4
O                 ATcT3EO   1    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] O <g> ATcT ver. 1.122, DHf298 = 249.229 � 0.002 kJ/mol - fit MAR17
 2.55160087E+00-3.83085457E-05 8.43197478E-10 4.01267136E-12-4.17476574E-16    2
 2.92287628E+04 4.87617014E+00 3.15906526E+00-3.21509999E-03 6.49255543E-06    3
-5.98755115E-09 2.06876117E-12 2.91298453E+04 2.09078344E+00 2.99753606E+04    4
!H                       H   1               G    300.00   4000.00 1000.00      1
! .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
! .254736600E+05-.446682850E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
! .000000000E+00 .000000000E+00 .254736600E+05-.446682850E+00                   4
H                 ATcT3EH   1    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] H <g> ATcT ver. 1.122, DHf298 = 217.998 � 0.000 kJ/mol - fit MAR17
 2.49985211E+00 2.34582548E-07-1.16171641E-10 2.25708298E-14-1.52992005E-18    2
 2.54738024E+04-4.45864645E-01 2.49975925E+00 6.73824499E-07 1.11807261E-09    3
-3.70192126E-12 2.14233822E-15 2.54737665E+04-4.45574009E-01 2.62191345E+04    4
!OH                      H   1O   1          G    300.00   4000.00 1000.00      1
! .283853033E+01 .110741289E-02-.294000209E-06 .420698729E-10-.242289890E-14    2
! .369780808E+04 .584494652E+01 .399198424E+01-.240106655E-02 .461664033E-05    3
!-.387916306E-08 .136319502E-11 .336889836E+04-.103998477E+00                   4
OH                ATcT3EH   1O   1    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] OH <g> ATcT ver. 1.122, DHf298 = 37.490 � 0.027 kJ/mol - fit MAR17
 2.84581721E+00 1.09723818E-03-2.89121101E-07 4.09099910E-11-2.31382258E-15    2
 3.71706610E+03 5.80339915E+00 3.97585165E+00-2.28555291E-03 4.33442882E-06    3
-3.59926640E-09 1.26706930E-12 3.39341137E+03-3.55397262E-02 4.50901087E+03    4
!HO2                     H   1O   2          G    300.00   4000.00 1000.00      1
! .417228741E+01 .188117627E-02-.346277286E-06 .194657549E-10 .176256905E-15    2
! .310206839E+02 .295767672E+01 .430179807E+01-.474912097E-02 .211582905E-04    3
!-.242763914E-07 .929225225E-11 .264018485E+03 .371666220E+01                   4
HO2               ATcT3EH   1O   2    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] HO2 <g> ATcT ver. 1.122, DHf298 = 12.26 � 0.16 kJ/mol - fit MAR17 
 4.10564010E+00 2.04046836E-03-3.65877562E-07 1.85973044E-11 4.98818315E-16    2
 4.32898769E+01 3.30808126E+00 4.26251250E+00-4.45642032E-03 2.05164934E-05    3
-2.35794011E-08 9.05614257E-12 2.62442356E+02 3.88223684E+00 1.47417835E+03    4
! C                       C   1               G    300.00   4000.00 1000.00      1
! .843301655E+00-.481886660E-02 .103261427E-04-.515161356E-08 .759963466E-12    2
! .868941443E+05 .170134676E+02 .000000000E+00 .000000000E+00 .000000000E+00    3
! .468280808E-08-.275232998E-11 .870122065E+05 .207811260E+02                   4
CSOLID                  C   1               G    300.00   4000.00 1000.00      1
 .159828070E+01 .143065097E-02-.509435105E-06 .864401302E-10-.534349530E-14    2
-.745940284E+03-.930332005E+01-.303744539E+00 .436036227E-02 .198268825E-05    3
-.643472598E-08 .299601320E-11-.109458288E+03 .108301475E+01                   4
CH                      C   1H   1          G    300.00   4000.00 1000.00      1
 .252093690E+01 .176536390E-02-.461476600E-06 .592896750E-10-.334745010E-14    2
 .709948780E+05 .740518290E+01 .348975830E+01 .324321600E-03-.168997510E-05    3
 .316284200E-08-.140618030E-11 .706607550E+05 .208428410E+01                   4
!HCO                     C   1H   1O   1     G    300.00   4000.00 1000.00      1
! .392001542E+01 .252279324E-02-.671004164E-06 .105615948E-09-.743798261E-14    2
! .365342928E+04 .358077056E+01 .423754610E+01-.332075257E-02 .140030264E-04    3
!-.134239995E-07 .437416208E-11 .387241185E+04 .330834869E+01                   4
HCO               ATcT3EC   1H   1O   1    0G    200.00   6000.00 1000.00      1	! [Ghobad] HCO <g> ATcT ver. 1.122, DHf298 = 41.803 � 0.099 kJ/mol - fit MAR17
 3.85781113E+00 2.64113950E-03-7.44177294E-07 1.23313230E-10-8.88958718E-15    2
 3.61642883E+03 3.92451197E+00 3.97074749E+00-1.49121608E-03 9.54041776E-06    3
-8.82720349E-09 2.67645129E-12 3.84203291E+03 4.44660361E+00 5.02774557E+03    4
HCO3                    C   1H   1O   3     G    300.00   4000.00 1000.00      1
 .726425669E+01 .532196974E-02-.196520055E-05 .323182996E-09-.195989250E-13    2
-.159242239E+05-.103647520E+02 .364808935E+01 .957717212E-02 .755287366E-05    3
-.181264650E-07 .827293980E-11-.146544449E+05 .967735548E+01                   4
CH2                     C   1H   2          G    300.00   4000.00 1000.00      1
 .314631886E+01 .303671259E-02-.996474439E-06 .150483580E-09-.857335515E-14    2
 .460412605E+05 .472341711E+01 .371757846E+01 .127391260E-02 .217347251E-05    3
-.348858500E-08 .165208866E-11 .458723866E+05 .175297945E+01                   4
CH2(S)                  C   1H   2          G    300.00   4000.00 1000.00      1
 .313501686E+01 .289593926E-02-.816668090E-06 .113572697E-09-.636262835E-14    2
 .505040504E+05 .406030621E+01 .419331325E+01-.233105184E-02 .815676451E-05    3
-.662985981E-08 .193233199E-11 .503662246E+05-.746734310E+00                   4
CH3                     C   1H   3          G    300.00   4000.00 1000.00      1
 .297812060E+01 .579785200E-02-.197558000E-05 .307297900E-09-.179174160E-13    2
 .165095130E+05 .472247990E+01 .365717970E+01 .212659790E-02 .545838830E-05    3
-.661810030E-08 .246570740E-11 .164227160E+05 .167353540E+01                   4
CH3O                    C   1H   3O   1     G    300.00   4000.00 1000.00      1
 .475779238E+01 .744142474E-02-.269705176E-05 .438090504E-09-.263537098E-13    2
 .390139164E+03-.196680028E+01 .371180502E+01-.280463306E-02 .376550971E-04    3
-.473072089E-07 .186588420E-10 .130772484E+04 .657240864E+01                   4
CH2OH                   C   1H   3O   1     G    300.00   4000.00 1000.00      1
 .509312037E+01 .594758550E-02-.206496524E-05 .323006703E-09-.188125052E-13    2
-.405813228E+04-.184690613E+01 .447832317E+01-.135069687E-02 .278483707E-04    3
-.364867397E-07 .147906775E-10-.352476728E+04 .330911984E+01                   4
CH3O2                   C   1H   3O   2     G    300.00   4000.00 1000.00      1
 .480390863E+01 .995844638E-02-.385301026E-05 .684740497E-09-.458402955E-13    2
-.747135460E+03 .145281400E+01 .362497097E+01 .359397933E-02 .226538097E-04    3
-.295391947E-07 .111977570E-10 .793040410E+02 .996382194E+01                   4
C2H                     C   2H   1          G    300.00   4000.00 1000.00      1
 .366270248E+01 .382492252E-02-.136632500E-05 .213455040E-09-.123216848E-13    2
 .671683790E+05 .392205792E+01 .289867676E+01 .132988489E-01-.280733327E-04    3
 .289484755E-07-.107502351E-10 .670616050E+05 .618547632E+01                   4
HCCO                    C   2H   1O   1     G    300.00   4000.00 1000.00      1
 .591479333E+01 .371408730E-02-.130137010E-05 .206473345E-09-.121476759E-13    2
 .193596301E+05-.550567269E+01 .187607969E+01 .221205418E-01-.358869325E-04    3
 .305402541E-07-.101281069E-10 .201633840E+05 .136968290E+02                   4
C2H3                    C   2H   3          G    300.00   4000.00 1000.00      1
 .415026763E+01 .754021341E-02-.262997847E-05 .415974048E-09-.245407509E-13    2
 .338566380E+05 .172812235E+01 .336377642E+01 .265765722E-03 .279620704E-04    3
-.372986942E-07 .151590176E-10 .344749589E+05 .791510092E+01                   4
CH3CO                   C   2H   3O   1     G    300.00   4000.00 1000.00      1
 .531371650E+01 .917377930E-02-.332203860E-05 .539474560E-09-.324523680E-13    2
-.364504140E+04-.167575580E+01 .403587050E+01 .877294870E-03 .307100100E-04    3
-.392475650E-07 .152968690E-10-.268207380E+04 .786176820E+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   4000.00 1000.00      1
 .653928338E+01 .780238629E-02-.276413612E-05 .442098906E-09-.262954290E-13    2
-.118858659E+04-.872091393E+01 .279502600E+01 .101099472E-01 .161750645E-04    3
-.310303145E-07 .139436139E-10 .162944975E+03 .123646657E+02                   4
CH3CO2                  C   2H   3O   2     G    300.00   4000.00 1000.00      1
 .700171955E+01 .101977290E-01-.365621800E-05 .589475086E-09-.352561321E-13    2
-.226135780E+05-.905267669E+01 .475563598E+01 .780915313E-02 .162272935E-04    3
-.241210787E-07 .942644561E-11-.215157456E+05 .478096491E+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   4000.00 1000.00      1
 .102188027E+02 .888408630E-02-.222887620E-05 .166265570E-09 .000000000E+00    2
-.256023886E+05-.219354293E+02 .384065500E+01 .218595100E-01-.904528040E-05    3
 .385393800E-09 .000000000E+00-.234946000E+05 .124829900E+02                   4
C2H5                    C   2H   5          G    300.00   4000.00 1000.00      1
 .432195633E+01 .123930542E-01-.439680960E-05 .703519917E-09-.418435239E-13    2
 .121759475E+05 .171103809E+00 .424185905E+01-.356905235E-02 .482667202E-04    3
-.585401009E-07 .225804514E-10 .129690344E+05 .444703782E+01                   4
PC2H4OH                 C   2H   5O   1     G    300.00   4000.00 1000.00      1
 .701348674E+01 .120204391E-01-.421992012E-05 .670675981E-09-.397135273E-13    2
-.616161779E+04-.862052409E+01 .420954137E+01 .912964578E-02 .247462263E-04    3
-.392945764E-07 .166541312E-10-.491511371E+04 .830445413E+01                   4
CH3OCH2                 C   2H   5O   1     G    300.00   4000.00 1000.00      1
 .594067593E+01 .129906358E-01-.456921036E-05 .726888932E-09-.430599587E-13    2
-.258503562E+04-.452841964E+01 .453195381E+01 .781884271E-02 .194968539E-04    3
-.274538336E-07 .106521135E-10-.170629244E+04 .506122980E+01                   4
SC2H4OH                 C   2H   5O   1     G    300.00   4000.00 1000.00      1
 .635842302E+01 .124356276E-01-.433096839E-05 .684530381E-09-.403713238E-13    2
-.953018581E+04-.605106112E+01 .422283250E+01 .512174798E-02 .348386522E-04    3
-.491943637E-07 .201183723E-10-.835622088E+04 .801675700E+01                   4
C2H5O2                  C   2H   5O   2     G    300.00   4000.00 1000.00      1
 .888872432E+01 .135833179E-01-.491116949E-05 .792343362E-09-.473525704E-13    2
-.744107388E+04-.190789836E+02 .450099327E+01 .687965342E-02 .474143971E-04    3
-.692287127E-07 .287395324E-10-.539547911E+04 .791490068E+01                   4
C2H4O2H                 C   2H   5O   2     G    300.00   4000.00 1000.00      1
 .941379980E+01 .133542122E-01-.468067639E-05 .743230845E-09-.439824231E-13    2
 .198459602E+04-.224516643E+02 .507456388E+01 .132389561E-01 .253758646E-04    3
-.438089546E-07 .189061540E-10 .371063204E+04 .272289544E+01                   4
DME-OO                  C   2H   5O   3     G    300.00   4000.00 1359.00      1
 .120501213E+02 .123072703E-01-.435221905E-05 .690896352E-09-.407091104E-13    2
-.227977573E+05-.323415629E+02 .515628105E+01 .216783339E-01-.561847228E-05    3
-.192807296E-08 .859447044E-12-.196244836E+05 .725163812E+01                   4
DME-QOOH                C   2H   5O   3     G    300.00   4000.00 1367.00      1
 .140894827E+02 .105710448E-01-.375281006E-05 .597314407E-09-.352604582E-13    2
-.191406716E+05-.429268872E+02 .543520255E+01 .272005914E-01-.150210893E-04    3
 .370396290E-08-.309396378E-12-.157034464E+05 .495012674E+01                   4
C2-OOQOOH               C   2H   5O   4     G    300.00   4000.00 1387.00      1
 .145471032E+02 .123393823E-01-.427259469E-05 .668763337E-09-.390196721E-13    2
-.196338761E+05-.408784236E+02 .590031872E+01 .305658528E-01-.185905950E-04    3
 .567871605E-08-.702799577E-12-.163916571E+05 .633051038E+01                   4
DME-OOQOOH              C   2H   5O   5     G    300.00   4000.00 1382.00      1
 .146274659E+02 .163794767E-01-.563311171E-05 .877481381E-09-.510186598E-13    2
-.370029335E+05-.399555488E+02 .771229157E+01 .301140957E-01-.165996092E-04    3
 .533577253E-08-.842885930E-12-.341808026E+05-.165902348E+01                   4
C3H2                    C   3H   2          G    300.00   4000.00 1000.00      1             ! Modified 1712
 .667324762E+01 .557728845E-02-.199180164E-05 .320289156E-09-.191216272E-13    2
 .607571184E+05-.972894405E+01 .243417332E+01 .173013063E-01-.118294047E-04    3
 .102756396E-08 .162626314E-11 .619074892E+05 .121012230E+02                   4
C3H3                    C   3H   3          G    300.00   4000.00 1000.00      1
 .714221719E+01 .761902211E-02-.267460030E-05 .424914904E-09-.251475443E-13    2
 .395709594E+05-.125848690E+02 .135110873E+01 .327411291E-01-.473827407E-04    3
 .376310220E-07-.118541128E-10 .407679941E+05 .152058598E+02                   4
C3H5-A                  C   3H   5          G    300.00   4000.00 1000.00      1
 .674633155E+01 .131071760E-01-.460059113E-05 .731029510E-09-.432759674E-13    2
 .171151431E+05-.125248814E+02 .165533607E+01 .163688750E-01 .210544223E-04    3
-.424018394E-07 .192638759E-10 .189454047E+05 .161040987E+02                   4
C3H5-T                  C   3H   5          G    300.00   4000.00 1000.00      1
 .611018050E+01 .146733950E-01-.536768220E-05 .869049320E-09-.519320060E-13    2
 .255324420E+05-.835557120E+01 .255440330E+01 .109867980E-01 .301743050E-04    3
-.472535680E-07 .197710730E-10 .271502420E+05 .132075920E+02                   4
C3H5-S                  C   3H   5          G    300.00   4000.00 1000.00      1
 .605091412E+01 .134052084E-01-.473450586E-05 .755380897E-09-.448421084E-13    2
 .290860210E+05-.673692060E+01 .333277282E+01 .106102499E-01 .217559727E-04    3
-.347145235E-07 .144476835E-10 .303404530E+05 .978922358E+01                   4
C3H5O                   C   3H   5O   1     G    300.00   4000.00 1402.00      1
 .102638186E+02 .117609932E-01-.389837957E-05 .592650815E-09-.338867417E-13    2
 .725938472E+04-.275108651E+02 .824068673E+00 .346749909E-01-.251786795E-04    3
 .956781953E-08-.148085302E-11 .104203725E+05 .228283070E+02                   4
RALD3                   C   3H   5O   1     G    300.00   4000.00 1366.00      1
 .979372730E+01 .168079281E-01-.684815970E-05 .118460585E-08-.738195109E-13    2
-.875662870E+04-.294639062E+02 .667614768E+01 .261082031E-02 .280410577E-04    3
-.226802600E-07 .516442572E-11-.510504908E+04-.439698728E+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   4000.00 1000.00      1
 .754410697E+01 .143443222E-01-.508381081E-05 .813200521E-09-.483673315E-13    2
-.748672286E+04-.114792587E+02 .470187196E+01 .551653762E-02 .427505858E-04    3
-.594680816E-07 .240685378E-10-.592845491E+04 .712932590E+01                   4
C3H5OO                  C   3H   5O   2     G    300.00   4000.00 1375.00      1
 .120289627E+02 .126220050E-01-.443107280E-05 .699998849E-09-.411059161E-13    2
 .440592543E+04-.346276747E+02 .316765415E+01 .300862111E-01-.169786280E-04    3
 .462955698E-08-.501220245E-12 .789477349E+04 .142601307E+02                   4
RALD3OO                 C   3H   5O   3     G    300.00   4000.00 1375.00      1
 .168446948E+02 .108808472E-01-.388442566E-05 .620614245E-09-.367342997E-13    2
-.242215993E+05-.597283331E+02 .351827789E+01 .399638014E-01-.273701195E-04    3
 .894188675E-08-.112554087E-11-.194047940E+05 .125456874E+02                   4
QALD3OO                 C   3H   5O   3     G    300.00   4000.00 1387.00      1
 .165672086E+02 .109861375E-01-.388980958E-05 .618066089E-09-.364435558E-13    2
-.159737374E+05-.559457656E+02 .175858492E+01 .494637636E-01-.434833502E-04    3
 .195880861E-07-.355128051E-11-.111728737E+05 .222887088E+02                   4
ZALD3OO                 C   3H   5O   5     G    300.00   4000.00 1387.00      1
 .207806034E+02 .116953349E-01-.414531832E-05 .659225856E-09-.388964379E-13    2
-.355954399E+05-.753605279E+02 .563102793E+01 .452923139E-01-.313606807E-04    3
 .100926022E-07-.119108613E-11-.302385330E+05 .649991022E+01                   4
NC3H7                   C   3H   7          G    300.00   4000.00 1000.00      1
 .649636579E+01 .177337992E-01-.624898046E-05 .995389495E-09-.590199770E-13    2
 .885973885E+04-.856389710E+01 .408211458E+01 .523240341E-02 .513554466E-04    3
-.699343598E-07 .281819493E-10 .104074558E+05 .839534919E+01                   4
IC3H7                   C   3H   7          G    300.00   4000.00 1000.00      1
 .530597255E+01 .189854588E-01-.674315384E-05 .107993730E-08-.642785036E-13    2
 .778748910E+04-.223233935E+01 .547421257E+01-.842536682E-02 .804607759E-04    3
-.949287824E-07 .359830971E-10 .904939013E+04 .340542323E+01                   4
CH3CH2CHOH              C   3H   7O   1     G   300.000  5000.000 1388.000    31 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
 1.14795375E+01 1.45881429E-02-4.88359380E-06 7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01 1.13614529E+00 3.68850655E-02-2.24073579E-05    3
 6.62398992E-09-7.32206246E-13-1.09273174E+04 2.24919343E+01                   4
CH3CH2CH2O              C   3H   7O   1    0G   300.000  5000.000 1386.000    21 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
 1.15279177E+01 1.53775991E-02-5.23946272E-06 8.11382512E-10-4.69927603E-14    2
-9.85099866E+03-3.54233008E+01 2.57486880E+00 3.07100600E-02-1.20048836E-05    3
 3.40807021E-12 7.25275283E-13-6.20913350E+03 1.45966401E+01                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   4000.00 1388.00      1
 .110944203E+02 .153549108E-01-.523574640E-05 .810964124E-09-.469665855E-13    2
-.134769536E+05-.307070215E+02 .584672920E+00 .407370189E-01-.294865043E-04    3
 .116950656E-07-.196228356E-11-.984929391E+04 .255429190E+02                   4
CH2CH2CH2OH             C   3H   7O   1    0G   300.000  5000.000 1402.000    31 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
 1.08178935E+01 1.53027604E-02-5.15746733E-06 7.92717531E-10-4.56680640E-14    2
-1.14319965E+04-2.79700973E+01 2.58072848E-01 3.90347698E-02-2.51378459E-05    3
 8.26896578E-09-1.09178202E-12-7.68516846E+03 2.90500173E+01                   4
CH3COHCH3               C   3H   7O   1     G    300.00   4000.00 1388.00      1
 .115026438E+02 .149881248E-01-.510421075E-05 .789864272E-09-.457135659E-13    2
-.164821894E+05-.347655748E+02 .118802517E+01 .410410262E-01-.314650841E-04    3
 .133514692E-07-.237788249E-11-.130177234E+05 .200655998E+02                   4
CH3CHCH2OH              C   3H   7O   1     G   300.000  5000.000 1393.000    31 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
 1.04922579E+01 1.55907665E-02-5.25786983E-06 8.08382729E-10-4.65762492E-14    2
-1.20531154E+04-2.64451618E+01 2.48398386E+00 3.14461742E-02-1.62613388E-05    3
 3.80532805E-09-2.66318786E-13-8.95721842E+03 1.76242658E+01                   4
NC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1374.00      1
 .146139980E+02 .143723015E-01-.488635144E-05 .756519620E-09-.438364992E-13    2
-.646101457E+04-.457478245E+02 .191005011E+01 .411666833E-01-.251630217E-04    3
 .711856873E-08-.698838732E-12-.179305093E+04 .234514457E+02                   4
IC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1399.00      1
 .155030898E+02 .139802008E-01-.481811216E-05 .751835399E-09-.437743118E-13    2
-.741643030E+04-.523911482E+02-.184042862E+00 .564670638E-01-.501611253E-04    3
 .230526863E-07-.423866481E-11-.252333896E+04 .298354826E+02                   4
NC3H7O2                 C   3H   7O   2     G    300.00   4000.00 1388.00      1
 .127230991E+02 .167336808E-01-.575943184E-05 .897769493E-09-.522275065E-13    2
-.108816595E+05-.381965321E+02 .156301709E+01 .426192697E-01-.296615075E-04    3
 .114187326E-07-.189894471E-11-.688086375E+04 .219842933E+02                   4
IC3H7O2                 C   3H   7O   2     G    300.00   4000.00 1392.00      1
 .132610651E+02 .162501084E-01-.558631798E-05 .870057473E-09-.505849469E-13    2
-.131937089E+05-.421023499E+02 .103495454E+01 .469942369E-01-.366525520E-04    3
 .157084173E-07-.281956117E-11-.906344820E+04 .229566921E+02                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1388.00      1
 .185146106E+02 .164157074E-01-.573085844E-05 .901975314E-09-.528299084E-13    2
-.231819444E+05-.618247164E+02 .254387733E+01 .570847379E-01-.472164204E-04    3
 .208289492E-07-.378162942E-11-.178600410E+05 .229447574E+02                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1391.00      1
 .191234208E+02 .158457151E-01-.552231946E-05 .868162288E-09-.508094203E-13    2
-.255253957E+05-.661419362E+02 .175906535E+01 .624712381E-01-.554930416E-04    3
 .257973727E-07-.483190839E-11-.200009572E+05 .251348546E+02                   4
C4H3                    C   4H   3          G    300.00   4000.00 1000.00      1
 .107527376E+02 .538115300E-02-.554963720E-06-.305226590E-09 .576173970E-13    2
 .612141980E+05-.297302533E+02 .415388100E+01 .172628700E-01-.238937390E-06    3
-.101870000E-07 .434050410E-11 .633807200E+05 .603650600E+01                   4
C4H3O                   C   4H   3O   1     G    300.00   4000.00 1000.00      1
 .129455763E+02 .795235476E-02-.280679691E-05 .445205248E-09-.262240810E-13    2
 .175946397E+05-.478819894E+02-.584674088E+01 .620875882E-01-.630010605E-04    3
 .306882361E-07-.575456234E-11 .230253176E+05 .492940922E+02                   4
C4H5                    C   4H   5          G    300.00   4000.00 1000.00      1
 .128659744E+02 .794336940E-02-.862646570E-06-.465563500E-09 .895113110E-13    2
 .378355213E+05-.418250446E+02 .299524000E+01 .228845610E-01 .197547090E-05    3
-.114824500E-07 .319782310E-11 .414221800E+05 .128945400E+02                   4
C4H71-4                 C   4H   7          G    300.00   4000.00 1000.00      1
 .664945270E+01 .226232110E-01-.806420670E-05 .954149200E-09 .000000000E+00    2
 .206794519E+05-.786429084E+01 .283048200E+00 .386777000E-01-.210739710E-04    3
 .427582900E-08 .000000000E+00 .225247800E+05 .254564400E+02                   4
IC4H7                   C   4H   7          G    300.00   4000.00 1000.00      1
 .616543300E+01 .257842760E-01-.936521250E-05 .112618500E-08 .000000000E+00    2
 .114713700E+05-.676561500E+01 .476952000E+01 .167724920E-01 .213011010E-04    3
-.275874430E-07 .845501100E-11 .126384700E+05 .401309300E+01                   4
C4H71-3                 C   4H   7          G    300.00   4000.00 1000.00      1
 .714879043E+01 .219663880E-01-.774471300E-05 .907477370E-09 .000000000E+00    2
 .124589843E+05-.117547735E+02-.442598200E+00 .422160100E-01-.254697900E-04    3
 .597432100E-08 .000000000E+00 .145672100E+05 .276086500E+02                   4
RALD4X                  C   4H   7O   1     G    300.00   4000.00 1378.00      1
 .109543855E+02 .241148701E-01-.952821930E-05 .161222652E-08-.988398314E-13    2
-.118963413E+05-.334390867E+02 .575601777E+01 .186084099E-01 .131646529E-04    3
-.151687447E-07 .367436225E-11-.792068905E+04 .141446613E+01                   4
RIBALDB                 C   4H   7O   1     G    300.00   4000.00 1000.00      1
 .355152000E+01 .294219200E-01-.104255000E-04 .171367900E-08-.107873000E-12    2
 .000000000E+00 .104367300E+02-.823550500E+00 .485680000E-01-.340648100E-04    3
 .109786600E-07-.495457100E-12 .000000000E+00 .303407900E+02                   4
RIBALDG                 C   4H   7O   1     G    300.00   4000.00 1000.00      1
 .499900800E+01 .269364000E-01-.923615800E-05 .148292200E-08-.918125000E-13    2
-.348819900E+04 .571944000E+01-.277712900E+01 .617368400E-01-.610123800E-04    3
 .338144900E-07-.767826900E-11-.241914600E+04 .416421800E+02                   4
RMP3                    C   4H   7O   2     G    300.00   4000.00 1376.00      1
 .154260382E+02 .169789201E-01-.593961909E-05 .936106835E-09-.548809672E-13    2
-.343012110E+05-.525677530E+02 .406577480E+01 .388324925E-01-.208048750E-04    3
 .506251249E-08-.421741752E-12-.297848227E+05 .102796868E+02                   4
QA4X                    C   4H   7O   3     G    300.00   4000.00 1000.00      1
 .778775690E+01 .301204420E-01-.104582260E-04 .169501670E-08-.105681860E-12    2
-.162963980E+05 .404129030E+00 .111242760E+01 .661709530E-01-.649819340E-04    3
 .331132210E-07-.636964220E-11-.160735140E+05 .288202740E+02                   4
RIBALDGOO               C   4H   7O   3     G    300.00   4000.00 1000.00      1
 .688742900E+01 .315358900E-01-.111087400E-04 .181743800E-08-.113981500E-12    2
-.209771000E+05 .101528900E+01-.131763500E+01 .654173000E-01-.523002100E-04    3
 .187106700E-07-.151244600E-11-.199258600E+05 .391267300E+02                   4
QIBALDB3                C   4H   7O   3     G    300.00   4000.00 1000.00      1
 0.77877569E+01 0.30120442E-01-0.10458226E-04 0.16950167E-08-0.10568186E-12    2
-0.16296398E+05 0.40412903E+00 0.11124276E+01 0.66170953E-01-0.64981934E-04    3
 0.33113221E-07-0.63696422E-11-0.16073514E+05 0.28820274E+02                   4
RIBALDBOO               C   4H   7O   3     G    300.00   4000.00 1000.00      1
 0.72319469E+01 0.32013219E-01-0.11485144E-04 0.19037878E-08-0.12050984E-12    2
-0.22166488E+05-0.72145844E+00-0.23625577E-01 0.64917222E-01-0.53189186E-04    3
 0.19445174E-07-0.16272577E-11-0.21545568E+05 0.31875837E+02                   4
QIBALDG3                C   4H   7O   3     G    300.00   4000.00 1000.00      1
 .815273500E+01 .289866500E-01-.985444500E-05 .157305600E-08-.970256900E-13    2
-.143742500E+05-.200325000E+01-.862350600E+00 .706020100E-01-.697863100E-04    3
 .360017200E-07-.720299500E-11-.133755300E+05 .389215900E+02                   4
QIBALDG2                C   4H   7O   3     G    300.00   4000.00 1000.00      1
 0.45559053E+01 0.35916157E-01-0.13290762E-04 0.22510276E-08-0.14461383E-12    2
-0.18124246E+05 0.16529331E+02 0.15762151E+01 0.67029655E-01-0.68767891E-04    3
 0.36980971E-07-0.75502798E-11-0.19410281E+05 0.24012136E+02                   4
RALD4OOX                C   4H   7O   3     G    300.00   4000.00 1000.00      1
 .723194690E+01 .320132190E-01-.114851440E-04 .190378780E-08-.120509840E-12    2
-.221664880E+05-.721458440E+00-.236255770E-01 .649172220E-01-.531891860E-04    3
 .194451740E-07-.162725770E-11-.215455680E+05 .318758370E+02                   4
ZIBALDB3                C   4H   7O   5     G    300.00   4000.00 1000.00      1
 .101088800E+02 .334733300E-01-.116762600E-04 .189872800E-08-.118662800E-12    2
-.318892400E+05-.778537800E+01 .612429000E+00 .741854800E-01-.608675100E-04    3
 .207212300E-07-.985714500E-12-.308839900E+05 .356398800E+02                   4
ZIBALDG2                C   4H   7O   5     G    300.00   4000.00 1000.00      1
 0.67585382E+01 0.40589843E-01-0.15337158E-04 0.26372311E-08-0.17129352E-12    2
-0.34054738E+05 0.10674515E+02 0.13726847E+01 0.78338057E-01-0.69229740E-04    3
 0.25735014E-07-0.17713571E-11-0.35033230E+05 0.29777508E+02                   4
ZA4X                    C   4H   7O   5     G    300.00   4000.00 1000.00      1
 .675853820E+01 .405898430E-01-.153371580E-04 .263723110E-08-.171293520E-12    2
-.340547380E+05 .106745150E+02 .137268470E+01 .783380570E-01-.692297400E-04    3
 .257350140E-07-.177135710E-11-.350332300E+05 .297775080E+02                   4
ZIBALDG3                C   4H   7O   5     G    300.00   4000.00 1000.00      1
 .101088800E+02 .334733300E-01-.116762600E-04 .189872800E-08-.118662800E-12    2
-.318892400E+05-.778537800E+01 .612429000E+00 .741854800E-01-.608675100E-04    3
 .207212300E-07-.985714500E-12-.308839900E+05 .356398800E+02                   4
PC4H9                   C   4H   9          G    300.00   4000.00 1000.00      1
 .285927140E+01 .339093470E-01-.129634890E-04 .162487360E-08 .000000000E+00    2
 .644131902E+04 .136765387E+02 .361027200E+00 .446560900E-01-.269622400E-04    3
 .737512580E-08 .000000000E+00 .679487900E+04 .252696800E+02                   4
TC4H9                   C   4H   9          G    300.00   4000.00 1000.00      1
 .678309830E+01 .275756420E-01-.999251920E-05 .119923980E-08 .000000000E+00    2
 .130943964E+04-.110379681E+02-.668177200E+00 .478197410E-01-.281268890E-04    3
 .654078610E-08 .000000000E+00 .334806900E+04 .274761900E+02                   4
SC4H9                   C   4H   9          G    300.00   4000.00 1000.00      1
 .182440000E+01 .354350280E-01-.136901980E-04 .172985780E-08 .000000000E+00    2
 .521137543E+04 .190721830E+02 .882678800E+00 .419813690E-01-.239577090E-04    3
 .639274900E-08 .000000000E+00 .513670700E+04 .226104800E+02                   4
IC4H9                   C   4H   9          G    300.00   4000.00 1000.00      1
 .672898190E+01 .277240280E-01-.100574610E-04 .120817530E-08 .000000000E+00    2
 .390175463E+04-.921990655E+01-.514098700E+00 .469939600E-01-.268680800E-04    3
 .599194290E-08 .000000000E+00 .591746700E+04 .283543100E+02                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   4000.00 1390.00      1
 .147487308E+02 .193476286E-01-.668165997E-05 .104395798E-08-.608330722E-13    2
-.178485397E+05-.492109234E+02 .467890397E+00 .521732276E-01-.362067190E-04    3
 .135025449E-07-.213961182E-11-.127480216E+05 .278224820E+02                   4
CH3CHCH2OCH3            C   4H   9O   1     G    300.00   4000.00 1422.00      1
 .148239632E+02 .195938055E-01-.674334212E-05 .105133556E-08-.611769464E-13    2
-.154937986E+05-.535942326E+02-.581327100E+00 .539666459E-01-.358338761E-04    3
 .122179671E-07-.171024843E-11-.995421675E+04 .297619860E+02                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   4000.00 1390.00      1
 .151619233E+02 .189741815E-01-.654734215E-05 .102237774E-08-.595503510E-13    2
-.208549516E+05-.532957109E+02 .108860217E+01 .524153990E-01-.380997951E-04    3
 .151074363E-07-.254404184E-11-.159195374E+05 .222613243E+02                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   4000.00 1422.00      1
 .140854789E+02 .197806925E-01-.671026390E-05 .103599950E-08-.598718336E-13    2
-.165129917E+05-.457671006E+02-.566170728E-01 .523981203E-01-.356379876E-04    3
 .128198684E-07-.192264202E-11-.115334457E+05 .303769293E+02                   4
CH3CH2CHCH2OH           C   4H   9O   1    0G   300.000  5000.000 1394.000    41 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 12_08_2016_14_12_47
+1.38348463E+01+1.99255957E-02-6.74388288E-06+1.03943751E-09-5.99954849E-14    2
-1.62408295E+04-4.28940661E+01+2.16591909E+00+4.43770980E-02-2.54941588E-05    3
+7.22842042E-09-7.87011274E-13-1.18784302E+04+2.08188392E+01+0.00000000E+00    4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   4000.00 1387.00      1
 .142049192E+02 .195897318E-01-.671801693E-05 .104483881E-08-.606940644E-13    2
-.190416934E+05-.463876157E+02 .933300006E+00 .472805232E-01-.278316313E-04    3
 .797039080E-08-.870532264E-12-.140666468E+05 .261224696E+02                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   4000.00 1390.00      1
 .147487308E+02 .193476286E-01-.668165997E-05 .104395798E-08-.608330722E-13    2
-.178485397E+05-.492109234E+02 .467890397E+00 .521732276E-01-.362067190E-04    3
 .135025449E-07-.213961182E-11-.127480216E+05 .278224820E+02                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   4000.00 1682.00      1
 .125605997E+02 .210637488E-01-.715019648E-05 .110439262E-08-.638428695E-13    2
-.183183621E+05-.368996627E+02 .329612707E+01 .347649647E-01-.102505618E-04    3
-.204641931E-08 .118879408E-11-.142607619E+05 .157499123E+02                   4
RTC4H8OH                C   4H   9O   1     G    300.00   4000.00 1395.00      1
 .146782533E+02 .193935063E-01-.660052048E-05 .102120044E-08-.590998119E-13    2
-.199408575E+05-.505292168E+02-.836665970E-01 .558040633E-01-.420184309E-04    3
 .171111519E-07-.290735214E-11-.149499995E+05 .281627857E+02                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   4000.00 1673.00      1
 .145354872E+02 .193544788E-01-.655352544E-05 .101052180E-08-.583473661E-13    2
-.195307842E+05-.500528678E+02 .524328525E+00 .528985884E-01-.379651080E-04    3
 .147054933E-07-.239054621E-11-.147012758E+05 .249822692E+02                   4
RTC4H9O                 C   4H   9O   1     G    300.00   4000.00 1391.00      1
 .154820006E+02 .191120896E-01-.659337031E-05 .102954283E-08-.599712426E-13    2
-.189474281E+05-.587209701E+02-.652960434E+00 .575360662E-01-.423660204E-04    3
 .165461682E-07-.269335532E-11-.133634774E+05 .277645681E+02                   4
CH3CH2CH2CHOH           C   4H   9O   1    0G   300.000  5000.000 1392.000    41 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 12_08_2016_14_12_47
+1.47813217E+01+1.89692972E-02-6.38671427E-06+9.81341181E-10-5.65332084E-14    2
-1.88487062E+04-4.98892364E+01+7.72566993E-01+5.00429367E-02-3.20163534E-05    3
+1.02913291E-08-1.30709217E-12-1.38421800E+04+2.58928300E+01+0.00000000E+00    4
CH3CH2CH2CH2O           C   4H   9O   1    0G   300.000  5000.000 1382.000    41 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 12_08_2016_14_12_47
+1.52662649E+01+1.94024981E-02-6.71808947E-06+1.05163276E-09-6.13656485E-14    2
-1.43012793E+04-5.43382882E+01+1.93228064E+00+4.47128724E-02-2.24881300E-05    3
+4.12226630E-09+3.99342930E-14-9.07148053E+03+1.93703892E+01+0.00000000E+00    4
CH3CHCH2CH2OH           C   4H   9O   1    0G   300.000  5000.000 1521.000    41 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 12_08_2016_14_12_47
+1.36682761E+01+1.97440068E-02-6.61586418E-06+1.01311840E-09-5.82212400E-14    2
-1.70603748E+04-4.19313460E+01+9.12869135E-01+4.43138287E-02-2.14369517E-05    3
+3.12967216E-09+3.57475931E-13-1.22046904E+04+2.82635095E+01+0.00000000E+00    4
CH3CH2CHOCH3            C   4H   9O   1     G    300.00   4000.00 1382.00      1
 .157118766E+02 .189436692E-01-.663728010E-05 .104718616E-08-.614402720E-13    2
-.169625442E+05-.584079611E+02-.123566480E+00 .537328693E-01-.359804830E-04    3
 .125064763E-07-.182873667E-11-.111514942E+05 .275750096E+02                   4
CH2CH2CH2CH2OH          C   4H   9O   1    0G   300.000  5000.000 1401.000    41 !\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 12_08_2016_14_12_47
+1.41519859E+01+1.96439700E-02-6.64537615E-06+1.02402720E-09-5.91001981E-14    2
-1.56141213E+04-4.43658958E+01-6.95634721E-02+5.20263179E-02-3.44849029E-05    3
+1.17704221E-08-1.63047436E-12-1.06053581E+04+3.22854711E+01+0.00000000E+00    4
IC4H9P-OO               C   4H   9O   2     G    300.00   4000.00 1391.00      1
 .160321835E+02 .211162441E-01-.726598082E-05 .113244436E-08-.658740064E-13    2
-.161760498E+05-.559920048E+02 .591660961E+00 .579744782E-01-.422019324E-04    3
 .167841571E-07-.283252682E-11-.107815683E+05 .268393730E+02                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   4000.00 1392.00      1
 .167547908E+02 .205266172E-01-.706765238E-05 .110199004E-08-.641203511E-13    2
-.197490954E+05-.625129056E+02 .429458545E+00 .619305024E-01-.492178248E-04    3
 .213391061E-07-.385156685E-11-.142778206E+05 .242205126E+02                   4
NC4H9-OO                C   4H   9O   2     G    300.00   4000.00 1392.00      1
 .164199470E+02 .207668293E-01-.714061871E-05 .111233445E-08-.646799300E-13    2
-.172909027E+05-.576444825E+02 .859225542E+00 .589774363E-01-.445935184E-04    3
 .184502497E-07-.321329944E-11-.119598721E+05 .254554544E+02                   4
NC4-QOOH                C   4H   9O   2     G    300.00   4000.00 1391.00      1
 .182943014E+02 .184250091E-01-.627217889E-05 .971379578E-09-.562825607E-13    2
-.128564704E+05-.650917535E+02 .986162058E+00 .585630676E-01-.416710545E-04    3
 .151223447E-07-.222454695E-11-.684048054E+04 .279289603E+02                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   4000.00 1396.00      1
 .181457399E+02 .188972595E-01-.650258715E-05 .101363925E-08-.589752496E-13    2
-.103249571E+05-.654833345E+02-.253900783E+00 .658110437E-01-.535280232E-04    3
 .228723790E-07-.398637599E-11-.429699727E+04 .319918975E+02                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   4000.00 1397.00      1
 .188631296E+02 .183239932E-01-.631233086E-05 .984688082E-09-.573186521E-13    2
-.138981290E+05-.708829284E+02-.425033602E+00 .698121411E-01-.606175877E-04    3
 .274812344E-07-.501908797E-11-.779203954E+04 .305104370E+02                   4
QBU1OOX                 C   4H   9O   3     G    300.00   4000.00 1386.00      1
 .129455763E+02 .795235476E-02-.280679691E-05 .445205248E-09-.262240810E-13    2
 .175946397E+05-.478819894E+02-.584674088E+01 .620875882E-01-.630010605E-04    3
 .306882361E-07-.575456234E-11 .230253176E+05 .492940922E+02                   4
RBU1OOX                 C   4H   9O   3     G    300.00   4000.00 1392.00      1
 .179101133E+02 .211247449E-01-.724787505E-05 .112742547E-08-.654930094E-13    2
-.371878276E+05-.612769774E+02 .289779336E+01 .560720331E-01-.390996379E-04    3
 .147174953E-07-.234862827E-11-.318812119E+05 .195265598E+02                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   4000.00 1391.00      1
 .225796674E+02 .201772761E-01-.702773819E-05 .110438266E-08-.646157968E-13    2
-.320684788E+05-.852469773E+02 .152317721E+01 .757827720E-01-.656981278E-04    3
 .300159936E-07-.556277284E-11-.252715176E+05 .257762885E+02                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   4000.00 1390.00      1
 .218612263E+02 .207812365E-01-.723484570E-05 .113659545E-08-.664871920E-13    2
-.284979533E+05-.798472350E+02 .156900216E+01 .724191880E-01-.596183448E-04    3
 .260680737E-07-.468228506E-11-.217597632E+05 .278260039E+02                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   4000.00 1393.00      1
 .231119306E+02 .196469811E-01-.682730172E-05 .107124796E-08-.626109519E-13    2
-.320261199E+05-.872192509E+02 .109604492E+01 .794472856E-01-.714221316E-04    3
 .334124791E-07-.626730135E-11-.251118713E+05 .282288973E+02                   4
ZBU1OOX                 C   4H   9O   5     G    300.00   4000.00 1397.00      1
 .236719411E+02 .205751255E-01-.708127339E-05 .110392970E-08-.642301320E-13    2
-.515463449E+05-.860806755E+02 .475209184E+01 .678608013E-01-.534336966E-04    3
 .221852722E-07-.378003417E-11-.452511232E+05 .144907043E+02                   4
C5H5                    C   5H   5          G    300.00   4000.00 1000.00      1
 .421464919E+01 .271834728E-01-.133173209E-04 .308980119E-08-.277879873E-12    2
 .288952416E+05-.305999781E-01-.737844042E+01 .972391818E-01-.169579138E-03    3
 .151818667E-06-.512075479E-10 .305514662E+05 .512829539E+02                   4
!C5H5O                   C   5H   5O   1     G    300.00   4000.00 1395.00      1       ! PROBABLY IT WAS 2,4 ISOMER. LEAST STABLE!!
! .149072105E+02 .136369619E-01-.470762207E-05 .736028654E-09-.429314124E-13    2
! .143724130E+05-.569296345E+02-.414628450E+01 .623584874E-01-.528374678E-04    3
! .224628793E-07-.380136191E-11 .204992627E+05 .437921058E+02                   4
C5H4OH Cyclo-2,4  T 5/10C  5.H  5.O  1.   0.G   200.000  6000.000 1000.        1
 1.32735713E+01 1.53094185E-02-5.50115205E-06 8.88634759E-10-5.32324947E-14    2
 2.27075873E+03-4.54766674E+01-1.74078500E+00 5.05423476E-02-1.59658908E-05    3
-2.73894335E-08 1.84710017E-11 6.52156699E+03 3.30332364E+01 8.06253742E+03    4
C5H4OH  Cyclo-2,4       H  5 C  5 O  1 N  0 G    200.0    3000.0   1000.0      1    ! DHof 20.16 LPM from automech C6H5+O2 paper
 8.15433468E+00 2.58109053E-02-1.32445071E-05 3.28780479E-09-3.19778186E-13    2
 4.12396691E+03-1.87762601E+01-3.76408182E-01 3.72784298E-02 1.39648368E-05    3
-5.42363862E-08 2.70582873E-11 6.75660088E+03 2.74100414E+01                   4
C5H4O                   H  4 C  5 O  1 N  0 G    200.0    3000.0   1000.0      1    ! DHof 16.41 LPM from automech C6H5+O2 paper
 6.54894513E+00 2.48908606E-02-1.27752734E-05 3.16512422E-09-3.06973283E-13    2
 3.28553663E+03-1.08667192E+01 6.45326515E-01 2.70140098E-02 2.70566468E-05    3
-6.20665862E-08 2.88732864E-11 5.32214959E+03 2.23237627E+01                   4
!C5H4OH Cyclo-2,4  T 5/10C  5.H  5.O  1.   0.G   200.000  6000.000 1000.        1 !burcat
! 1.32735713E+01 1.53094185E-02-5.50115205E-06 8.88634759E-10-5.32324947E-14    2
! 2.27075873E+03-4.54766674E+01-1.74078500E+00 5.05423476E-02-1.59658908E-05    3
!-2.73894335E-08 1.84710017E-11 6.52156699E+03 3.30332364E+01 8.06253742E+03    4
C5H5O  1-oxy-1,3- T09/10C  5.H  5.O  1.   0.G   200.000  6000.000 1000.        1
 1.14579913E+01 1.74857813E-02-6.31033387E-06 1.02222611E-09-6.13529798E-14    2
-7.47305910E+02-3.63570579E+01 1.02688782E+00 2.49799222E-02 4.13379251E-05    3
-7.92827590E-08 3.55323358E-11 3.01148270E+03 2.22500883E+01 4.65324451E+03    4
!C5H5O  1-oxy-1,4- T09/10C  5.H  5.O  1.   0.G   200.000  6000.000 1000.        1
! 1.14306204E+01 1.75353472E-02-6.33385273E-06 1.02662642E-09-6.16410846E-14    2
! 3.35973647E+03-3.62255087E+01 9.94952201E-01 2.57061151E-02 3.87827528E-05    3
!-7.61408558E-08 3.42541359E-11 7.09986737E+03 2.22760126E+01 8.74741530E+03    4
!C5H5O Cyclo-2,4-  T 3/10C  5.H  5.O  1.   0.G   200.000  6000.000 1000.        1      produced from C5H5+HO2
! 1.20244667E+01 1.69698914E-02-6.12274609E-06 9.91737990E-10-5.95206422E-14    2
! 2.05122293E+04-3.95370458E+01 7.74871946E-01 2.53185105E-02 4.65761215E-05    3
!-8.92691495E-08 4.04034749E-11 2.44938481E+04 2.34455624E+01 2.61043645E+04    4
C5H5OH Cyclo-1,3  T 8/10C  5.H  6.O  1.   0.G   200.000  6000.000 1000.        1
 1.20653902E+01 1.87856222E-02-6.69025883E-06 1.07435931E-09-6.40970640E-14    2
-1.02087893E+04-3.99330360E+01-4.45002464E-01 3.67965171E-02 2.13479506E-05    3
-6.30989227E-08 3.05704733E-11-6.13350745E+03 2.81881469E+01-4.55234957E+03    4
!C5H5OH Cyclo-1,4  T 8/10C  5.H  6.O  1.   0.G   200.000  6000.000 1000.        1
! 1.21107707E+01 1.87471485E-02-6.67696496E-06 1.07227634E-09-6.39751958E-14    2
!-1.06517616E+04-4.02092317E+01-6.03126120E-01 3.76204145E-02 2.01258044E-05    3
!-6.24427856E-08 3.04889481E-11-6.54057343E+03 2.88740619E+01-4.97947985E+03    4
!C5H5OH Cyclo-2,4  T 8/10C  5.H  6.O  1.   0.G   200.000  6000.000 1000.        1
! 1.16115218E+01 1.91901010E-02-6.83602335E-06 1.09795484E-09-6.55125692E-14    2
!-5.69452475E+03-3.68452441E+01 2.28105979E+00 1.72605889E-02 6.60492754E-05    3
!-1.06481809E-07 4.58889262E-11-1.99035320E+03 1.74654781E+01-1.48297975E+02    4
C5H7                    C   5H   7          G    300.00   4000.00 1000.00      1
 .671323690E+01 .274278890E-01-.994311090E-05 .119373240E-08 .000000000E+00    2
 .235116384E+05-.112735252E+02 .759315300E+00 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .251686000E+05 .196131100E+02                   4
RMCROTA                 C   5H   7O   2     G    300.00   4000.00 1000.00      1
 .151681730E+02 .178142000E-01-.496258460E-05 .688767770E-09-.386765100E-13    2
-.320532540E+05-.462913590E+02-.242828070E+00 .630479530E-01-.556979940E-04    3
 .265678430E-07-.501508770E-11-.278218120E+05 .329157640E+02                   4
NC5H9-3                 C   5H   9          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
ERC4H8CHO               C   5H   9O   1     G    300.00   4000.00 1517.00      1
 .190577032E+02 .197405268E-01-.706907553E-05 .113169306E-08-.670771090E-13    2
-.128899482E+05-.729817022E+02 .467212037E+01 .343554368E-01 .295219352E-05    3
-.145463894E-07 .444316435E-11-.603466621E+04 .109564879E+02                   4
C5EN-QOOH               C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OO                 C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
RMBX                    C   5H   9O   2     G    300.00   4000.00 1382.00      1
 .193382201E+02 .209401493E-01-.732209753E-05 .115371679E-08-.676297088E-13    2
-.412852468E+05-.755834444E+02 .231680806E+01 .569247905E-01-.356059275E-04    3
 .110212330E-07-.136558032E-11-.349304634E+05 .172843303E+02                   4
RMBOOX                  C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .211938570E+02 .222144000E-01-.631327380E-05 .888168590E-09-.502931100E-13    2
-.572489530E+05-.734085620E+02 .256566330E+01 .606897660E-01-.678613150E-05    3
-.390168040E-07 .205529000E-10-.518452190E+05 .251823650E+02                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
QMBOOX                  C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .211938570E+02 .222144000E-01-.631327380E-05 .888168590E-09-.502931100E-13    2
-.572489530E+05-.734085620E+02 .256566330E+01 .606897660E-01-.678613150E-05    3
-.390168040E-07 .205529000E-10-.518452190E+05 .251823650E+02                   4
ZMBOOX                  C   5H   9O   6     G    300.00   4000.00 1000.00      1
 .261471200E+02 .215283560E-01-.581135510E-05 .785452200E-09-.431572980E-13    2
-.689643590E+05-.913329620E+02 .443715430E+01 .699071290E-01-.165602940E-04    3
-.356586160E-07 .205531550E-10-.628690510E+05 .226288070E+02                   4
NC5H11                  C   5H  11          G    300.00   4000.00 1384.00      1
 .131340658E+02 .260923466E-01-.897731137E-05 .139920325E-08-.813970860E-13    2
-.427735231E+04-.434455998E+02-.304386354E+01 .581995422E-01-.316090839E-04    3
 .790004927E-08-.665198232E-12 .199185425E+04 .455946950E+02                   4
IC5H11                  C   5H  11          G    300.00   4000.00 1389.00      1
 .153818750E+02 .241141042E-01-.827847584E-05 .128831856E-08-.748649188E-13    2
-.184296128E+04-.564907641E+02-.592409395E+00 .586734947E-01-.365981110E-04    3
 .118412541E-07-.159845819E-11 .405970723E+04 .304115490E+02                   4
NEOC5H11                C   5H  11          G    300.00   4000.00 1396.00      1
 .166235914E+02 .227037884E-01-.771624835E-05 .119289853E-08-.690060600E-13    2
-.396429146E+04-.644693953E+02-.158140132E+01 .657175067E-01-.468120314E-04    3
 .174732793E-07-.268709925E-11 .230933742E+04 .331296742E+02                   4
RIPENTOHB               C   5H  11O   1     G    300.00   4000.00 1374.00      1
 .178146436E+02 .231777549E-01-.776038398E-05 .118900766E-08-.683934164E-13    2
-.225247765E+05-.648614694E+02 .204135308E+00 .588299650E-01-.324898705E-04    3
 .750026128E-08-.365893927E-12-.159312048E+05 .315479677E+02                   4
RIPENTOHA               C   5H  11O   1     G    300.00   4000.00 1394.00      1
 .176264597E+02 .239817014E-01-.815640882E-05 .126137771E-08-.729792490E-13    2
-.238094100E+05-.651182426E+02 .287733983E+00 .650700888E-01-.461663158E-04    3
 .176228098E-07-.282635934E-11-.177872581E+05 .278924962E+02                   4
RPENT1O                 C   5H  11O   1     G    300.00   5000.00 1396.00      1!\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
+1.87118024E+01+2.36054696E-02-8.05610528E-06+1.24900841E-09-7.23989034E-14    2
-1.84133036E+04-7.11769229E+01+1.61443159E+00+5.84449099E-02-3.26027513E-05    3
+7.76525028E-09-4.48739932E-13-1.20210227E+04+2.23620686E+01                   4
RPENT1OHB               C   5H  11O   1     G    300.00   5000.00 1394.00      1!\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
+1.71780951E+01+2.42601001E-02-8.22986526E-06+1.27049816E-09-7.34155598E-14    2
-2.04290445E+04-5.93472290E+01+1.84753679E+00+5.73086840E-02-3.47271444E-05    3
+1.06516139E-08-1.30777652E-12-1.47995754E+04+2.40150308E+01                   4
RPENT1OHE               C   5H  11O   1     G    300.00   5000.00 1400.00      1!\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
+1.74868543E+01+2.39842944E-02-8.13298324E-06+1.25529418E-09-7.25301446E-14    2
-1.97969015E+04-6.07667197E+01-3.94307020E-01+6.50012333E-02-4.38043364E-05    3
+1.52539819E-08-2.16516288E-12-1.35258816E+04+3.55083245E+01                   4
RPENT1OHD               C   5H  11O   1     G    300.00   5000.00 2022.00      1!\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
 1.65897836E+01 2.53826913E-02-9.43220215E-06 1.55249347E-09-9.39190299E-14    2
-2.10435752E+04-5.62532844E+01 3.69891615E-01 5.63524034E-02-2.76588983E-05    3
 4.35237097E-09 2.03539591E-13-1.50416080E+04 3.28904903E+01                   4
RIPENTO                 C   5H  11O   1     G    300.00   4000.00 1390.00      1
 .179852494E+02 .240897408E-01-.828641852E-05 .129144549E-08-.751291843E-13    2
-.197891737E+05-.690290731E+02-.769895465E+00 .660085470E-01-.438697957E-04    3
 .150115512E-07-.211319317E-11-.130499892E+05 .324309009E+02                   4
RPENT1OHA               C   5H  11O   1     G    300.00   5000.00 1394.00      1!\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
+1.80953018E+01+2.33361161E-02-7.88463541E-06+1.21428332E-09-7.00616136E-14    2
-2.30206675E+04-6.61675776E+01+4.26049539E-01+6.31258286E-02-4.15122762E-05    3
+1.38895665E-08-1.86732010E-12-1.67596661E+04+2.92144308E+01                   4
RIPENTOHD               C   5H  11O   1     G    300.00   4000.00 1394.00      1
 .172306012E+02 .242975217E-01-.826186089E-05 .127755536E-08-.739123165E-13    2
-.208013525E+05-.618034685E+02-.237764707E+00 .644135904E-01-.436552710E-04    3
 .156133960E-07-.232736806E-11-.146304196E+05 .323161057E+02                   4
RPENT1OHC               C   5H  11O   1     G    300.00   5000.00 1042.00      1!\AUTHOR: CR/KPS !\REF: GA !\COMMENT: FITTED WITH THERM ON 11_08_2016_20_43_11
+1.68143234E+01+2.44876194E-02-8.29372543E-06+1.27921101E-09-7.38804613E-14    2
-2.12567818E+04-5.74573295E+01+5.41167712E-01+5.66862244E-02-2.94678472E-05    3
+5.84904634E-09-3.31866470E-14-1.50943752E+04+3.18827465E+01                   4
RIPENTOHC               C   5H  11O   1     G    300.00   4000.00 1381.00      1
 .157053942E+02 .255921700E-01-.870811298E-05 .134716260E-08-.779628294E-13    2
-.226082350E+05-.522449991E+02 .309642922E+01 .468661615E-01-.183869508E-04    3
 .820832987E-09 .767460794E-12-.173551008E+05 .184684107E+02                   4
RMTBE                   C   5H  11O   1     G    300.00   4000.00 1386.00      1
 .191923401E+02 .226496418E-01-.770522799E-05 .119249279E-08-.690514122E-13    2
-.223486482E+05-.717004889E+02-.284403552E+00 .706092470E-01-.543641242E-04    3
 .224557925E-07-.385680161E-11-.157511970E+05 .321647207E+02                   4
NEOC5H11-OO             C   5H  11O   2     G    300.00   4000.00 1396.00      1
 .202154849E+02 .245786365E-01-.841704919E-05 .130775217E-08-.759095109E-13    2
-.224777899E+05-.796085899E+02 .730403748E+00 .705036948E-01-.502866599E-04    3
 .189083885E-07-.294948183E-11-.157211898E+05 .249439750E+02                   4
NEOC5-QOOH              C   5H  11O   2     G    300.00   4000.00 1396.00      1
 .218550366E+02 .228989820E-01-.786956915E-05 .122572909E-08-.712760383E-13    2
-.164801773E+05-.857429310E+02 .115441893E+01 .724266160E-01-.535668095E-04    3
 .205704339E-07-.323425526E-11-.941504872E+04 .250054329E+02                   4
NC5-QOOH                C   5H  11O   2     G    300.00   4000.00 1396.00      1
 .220245928E+02 .228314385E-01-.786198359E-05 .122609365E-08-.713571493E-13    2
-.179960313E+05-.864387261E+02-.607426660E+00 .818016374E-01-.685494236E-04    3
 .302071532E-07-.540750321E-11-.106868081E+05 .330450153E+02                   4
NC5H12OO                C   5H  11O   2     G    300.00   4000.00 1392.00      1
 .199150940E+02 .250390538E-01-.861981469E-05 .134386616E-08-.781893344E-13    2
-.238472344E+05-.769667628E+02 .235935841E+00 .739755736E-01-.572379508E-04    3
 .241234657E-07-.425357119E-11-.171710700E+05 .279024996E+02                   4
RPENT1OOX               C   5H  11O   3     G    300.00   4000.00 1394.00      1
 .235310388E+02 .257989924E-01-.888660144E-05 .138620388E-08-.806892959E-13    2
-.591984578E+05-.904223960E+02 .177546391E+01 .768095280E-01-.550828141E-04    3
 .206638345E-07-.320646569E-11-.516288295E+05 .264068764E+02                   4
QIPENTOOX               C   5H  11O   3     G    300.00   4000.00 1393.00      1
 .229723533E+02 .230366475E-01-.771154566E-05 .118147984E-08-.679624947E-13    2
-.349052726E+05-.847531774E+02 .275419521E+01 .666225847E-01-.414002404E-04    3
 .119392262E-07-.118354877E-11-.276318447E+05 .249380687E+02                   4
RIPENTOOX               C   5H  11O   3     G    300.00   4000.00 1394.00      1
 .229563234E+02 .264776592E-01-.906923239E-05 .140937564E-08-.818234063E-13    2
-.583968852E+05-.878789834E+02 .176378684E+01 .755411075E-01-.526303110E-04    3
 .191090062E-07-.286212429E-11-.509737373E+05 .261265484E+02                   4
MTBE-OO                 C   5H  11O   3     G    300.00   4000.00 1386.00      1
 .219476262E+02 .253064866E-01-.877948807E-05 .137597948E-08-.803553517E-13    2
-.383949561E+05-.811182382E+02 .226233362E+01 .712292692E-01-.511734982E-04    3
 .199100134E-07-.329751069E-11-.314029562E+05 .248780910E+02                   4
QPENT1OOX               C   5H  11O   3     G    300.00   4000.00 1393.00      1
 .246066807E+02 .226714906E-01-.788343040E-05 .123763348E-08-.723672450E-13    2
-.382649798E+05-.958452159E+02 .148247361E+01 .786233062E-01-.604614335E-04    3
 .240553703E-07-.391498689E-11-.304133501E+05 .276855455E+02                   4
MTBE-QOOH               C   5H  11O   3     G    300.00   4000.00 1401.00      1
 .214971173E+02 .259064341E-01-.848605930E-05 .127921441E-08-.726936886E-13    2
-.312441531E+05-.765479844E+02 .134883146E+01 .795292274E-01-.643595941E-04    3
 .280404405E-07-.497823206E-11-.249060790E+05 .293286141E+02                   4
NEOC5-OOQOOH            C   5H  11O   4     G    300.00   4000.00 1392.00      1
 .248490803E+02 .252599638E-01-.873651764E-05 .136662251E-08-.797082603E-13    2
-.350133010E+05-.961825156E+02 .265748524E+01 .758789336E-01-.526594216E-04    3
 .186692316E-07-.269820831E-11-.271776626E+05 .234450387E+02                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   4000.00 1391.00      1
 .257270270E+02 .247172056E-01-.859292907E-05 .134865114E-08-.788382618E-13    2
-.361631686E+05-.100728579E+03 .135798731E+01 .877212925E-01-.735867140E-04    3
 .327395450E-07-.595540146E-11-.281695250E+05 .282261555E+02                   4
ZIPENTOOX               C   5H  11O   5     G    300.00   4000.00 1400.00      1
 .258845592E+02 .261151092E-01-.903875069E-05 .141449719E-08-.825222954E-13    2
-.550208255E+05-.962071206E+02 .391413178E+01 .765170930E-01-.535251760E-04    3
 .194861484E-07-.294077918E-11-.472474207E+05 .222011325E+02                   4
MTBE-OOQOOH             C   5H  11O   5     G    300.00   4000.00 1391.00      1
 .264681284E+02 .261757287E-01-.899393547E-05 .140058534E-08-.814301239E-13    2
-.504985383E+05-.992053288E+02 .454595241E+01 .801871705E-01-.616423289E-04    3
 .254521416E-07-.437448229E-11-.430642384E+05 .177072264E+02                   4
ZPENT1OOX               C   5H  11O   5     G    300.00   4000.00 1400.00      1
 .286303066E+02 .232317088E-01-.801616025E-05 .125197153E-08-.729415409E-13    2
-.577713687E+05-.109745016E+03 .345682525E+01 .876757175E-01-.724014952E-04    3
 .308846552E-07-.532198779E-11-.496056070E+05 .234305819E+02                   4
C6H3                    C   6H   3          G    300.00   4000.00 1000.00      1
 .120132339E+02 .114461128E-01-.408884040E-05 .657753914E-09-.392832116E-13    2
 .825892145E+05-.335118700E+02 .150089155E+01 .545901804E-01-.788221454E-04    3
 .627969099E-07-.200768594E-10 .849133510E+05 .176237455E+02                   4
!C6H5                    C   6H   5          G    300.00   4000.00 1000.00      1 !polimi
! .157758892E+02 .965110900E-02-.942941600E-06-.546911100E-09 .102652200E-12    2
! .330269797E+05-.617628096E+02 .114355700E+00 .362732400E-01 .115828600E-05    3
!-.219696400E-07 .846355600E-11 .383605400E+05 .238011700E+02                   4
!C6H5 phenyl radi  T07/10C  6.H  5.   0.   0.G   200.000  6000.000  B  77.10390 1 
C6H5                    C   6H   5          G    300.00   4000.00 1000.00      1 !Burcat kik
 1.09540673E+01 1.82072569E-02-6.63331157E-06 1.08125690E-09-6.51736617E-14    2
 3.51098413E+04-3.64320659E+01 4.91024498E-01 1.72669813E-02 7.02556406E-05    3
-1.13389805E-07 4.89202543E-11 3.92340510E+04 2.42505364E+01 4.05676342E+04    4
LC6H5                   C   6H   5          G    300.00   4000.00 1000.00      1
 .134117680E+02 .147202210E-01-.508177050E-05 .798863540E-09-.469508440E-13    2
 .585037160E+05-.416520320E+02 .779297070E+00 .543721260E-01-.478738140E-04    3
 .161871640E-07 .337357440E-12 .616503120E+05 .221285920E+02                   4
C6H5O                   H   5C   6O   1     G   100.000  5000.000 1045.70      1 !UPDATED RDB - Currane
 1.13847939E+01 2.20913987E-02-9.35923352E-06 1.81143777E-09-1.31169823E-13    2
 1.06782097E+03-3.61613841E+01 2.03763899E+00 3.28240830E-02 1.11381131E-05    3
-3.41391653E-08 1.39344349E-11 4.39073906E+03 1.58922741E+01                   4
!C6H5O                   C   6H   5O   1     G    300.00   4000.00 1000.00      1
! .137221720E+02 .174688771E-01-.635504520E-05 .103492308E-08-.623410504E-13    2
! .287274751E+03-.488181680E+02-.466204455E+00 .413443975E-01 .132412991E-04    3
!-.572872769E-07 .289763707E-10 .477858391E+04 .276990274E+02                   4
DMF-3YL                 C   6H   7O   1     G    300.00   4000.00 1000.00      1
 .118002735E+02 .257930235E-01-.101089409E-04 .181299326E-08-.122176870E-12    2
 .130508362E+05-.352008048E+02 .197118616E+01 .384836786E-01 .786460722E-05    3
-.354301012E-07 .162325679E-10 .165648455E+05 .193223377E+02                   4
CYC6H9                  C   6H   9          G    300.00   4000.00 1381.00      1
 .166730638E+02 .227088190E-01-.801509353E-05 .127088484E-08-.748275111E-13    2
 .698387216E+04-.723601536E+02-.631908086E+01 .726795534E-01-.484456826E-04    3
 .157628084E-07-.202092558E-11 .153574632E+05 .524769640E+02                   4
RC6H9A                  C   6H   9          G    300.00   4000.00 1400.00      1
 .170842767E+02 .208842788E-01-.714529004E-05 .110943563E-08-.643676989E-13    2
 .201040204E+05-.639326012E+02-.266715213E+01 .726196475E-01-.605323920E-04    3
 .266000571E-07-.474613408E-11 .264415017E+05 .402220332E+02                   4
RALDEST                 C   6H   9O   3     G    300.00   4000.00 1373.00      1
 .215153215E+02 .236419666E-01-.830694270E-05 .131026314E-08-.767602984E-13    2
-.530993462E+05-.770487448E+02 .687062608E+01 .492844450E-01-.217786396E-04    3
 .243527207E-08 .464021620E-12-.470662293E+05 .479532953E+01                   4
CYC6H11                 C   6H  11          G    300.00   4000.00 1674.00      1
 .146799252E+02 .309324453E-01-.112934485E-04 .183887582E-08-.110464203E-12    2
-.197594614E+03-.590168221E+02-.757310296E+01 .766896480E-01-.424441426E-04    3
 .941423236E-08-.439999709E-12 .764576045E+04 .620172120E+02                   4
CYC6-QOOH-4             C   6H  11O   2     G    300.00   4000.00 1374.00      1
 .241250295E+02 .262273012E-01-.925328534E-05 .146724451E-08-.864028312E-13    2
-.163808524E+05-.106267870E+03-.596804450E+01 .893075551E-01-.558813589E-04    3
 .152003723E-07-.125762311E-11-.534935832E+04 .576800888E+02                   4
CYC6-OO                 C   6H  11O   2     G    300.00   4000.00 1380.00      1
 .225527144E+02 .280656231E-01-.990087442E-05 .156942170E-08-.923867180E-13    2
-.209455781E+05-.994788807E+02-.594021024E+01 .887171975E-01-.569424328E-04    3
 .171601250E-07-.191055830E-11-.104841379E+05 .556048484E+02                   4
CYC6-QOOH-2             C   6H  11O   2     G    300.00   4000.00 1375.00      1
 .243899542E+02 .262326944E-01-.930434909E-05 .148019558E-08-.873538395E-13    2
-.163135893E+05-.107549099E+03-.378907832E+01 .841562901E-01-.510965662E-04    3
 .133666762E-07-.102528616E-11-.580881865E+04 .464783226E+02                   4
CYC6-QOOH-3             C   6H  11O   2     G    300.00   4000.00 1374.00      1
 .241250295E+02 .262273012E-01-.925328534E-05 .146724451E-08-.864028312E-13    2
-.163808524E+05-.106267870E+03-.596804450E+01 .893075551E-01-.558813589E-04    3
 .152003723E-07-.125762311E-11-.534935832E+04 .576800888E+02                   4
CYC6-OOQOOH-4           C   6H  11O   4     G    300.00   4000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128893429E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .565320100E+02                   4
CYC6-OOQOOH-3           C   6H  11O   4     G    300.00   4000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128198915E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .572265244E+02                   4
CYC6-OOQOOH-2           C   6H  11O   4     G    300.00   4000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128198915E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .572265244E+02                   4
RDIPE                   C   6H  13O   1     G    300.00   4000.00 1389.00      1
 .195346832E+02 .300586517E-01-.103564671E-04 .161544621E-08-.940217507E-13    2
-.289625035E+05-.700231442E+02-.545711430E-01 .748436725E-01-.509801332E-04    3
 .191769721E-07-.313046382E-11-.218696353E+05 .358513387E+02                   4
!C7H7                    C   7H   7          G    300.00   4000.00 1000.00      1 ! Polimi
! .126890424E+02 .248754040E-01-.820402330E-05 .901804910E-09 .000000000E+00    2
! .179417186E+05-.454264236E+02-.296228400E+01 .659171040E-01-.433334430E-04    3
! .106408510E-07 .000000000E+00 .223472400E+05 .359657700E+02                   4
C7H7 Benzyl rad   T08/90C   7H   7    0    0G   200.000  6000.000 1000.        1 ! Burcat kik
 0.14043980E+02 0.23493873E-01-0.85375367E-05 0.13890841E-08-0.83614420E-13    2
 0.18564203E+05-0.51665589E+02 0.48111540E+00 0.38512832E-01 0.32861492E-04    3
-0.76972721E-07 0.35423068E-10 0.23307027E+05 0.23548820E+02 0.25317186E+05    4
!CH3C6H4                 C   7H   7          G    300.00   4000.00 1000.00      1 POLIMI
! .989521100E+01 .281997140E-01-.985390310E-05 .114532240E-08 .000000000E+00    2
! .307512908E+05-.257557742E+02-.298827000E+01 .621039310E-01-.390118950E-04    3
! .928257830E-08 .000000000E+00 .343676800E+05 .412025200E+02                   4
CH3C6H4 o-Tolu RadT10/13C  7.H  7.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat kik  1706
 1.28543060E+01 2.42712778E-02-8.75277064E-06 1.41703290E-09-8.50082345E-14    2
 3.10872386E+04-4.29177096E+01 2.43474215E+00 2.10368651E-02 7.20305506E-05    3
-1.14038924E-07 4.82416036E-11 3.53949018E+04 1.83045052E+01 3.74896416E+04    4
!
!CH3C6H4                 C   7H   7    0    0G   300.000  5000.000 1393.000    11      !Zhang
! 1.50088040E+01 2.08076711E-02-7.18274868E-06 1.12201995E-09-6.53756838E-14    2
! 2.89360689E+04-5.63866198E+01-2.51731357E+00 6.18263711E-02-4.43238513E-05    3
! 1.66517959E-08-2.59379321E-12 3.50509401E+04 3.77723973E+01                   4
!
OC6H4CH3                C   7H   7O   1     G    300.00   4000.00 1000.00      1
 .632623400E+01 .370920700E-01-.137369600E-04 .232847100E-08-.149701800E-12    2
-.156635900E+04-.468621100E+01-.403964400E+01 .739909500E-01-.515945300E-04    3
 .120372800E-07 .143210200E-11 .225707600E+03 .453169300E+02                   4
HOC6H4CH2               C   7H   7O   1     G    300.00   4000.00 1000.00      1
 .689970000E+01 .376640500E-01-.142499000E-04 .245139600E-08-.159215300E-12    2
-.104378100E+04-.796692700E+01-.415304900E+01 .776998800E-01-.583028700E-04    3
 .178677900E-07-.536299700E-12 .896696700E+03 .453288900E+02                   4
RMCYC6                  C   7H  13          G    300.00   4000.00 2030.00      1
 .173202469E+02 .361144629E-01-.130438584E-04 .210911191E-08-.126098895E-12    2
-.514813032E+04-.717714814E+02-.853970231E+01 .919151844E-01-.546389770E-04    3
 .144889205E-07-.127842414E-11 .374687760E+04 .679730355E+02                   4
NC7H13                  C   7H  13          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
MCYC6-QOOH              C   7H  13O   2     G    300.00   4000.00 2055.00      1
 .234331685E+02 .347621964E-01-.124048044E-04 .199225952E-08-.118633947E-12    2
-.195868561E+05-.990888361E+02-.694095755E+01 .104651350E+00-.698281467E-04    3
 .219897276E-07-.260222584E-11-.958151058E+04 .634587763E+02                   4
RMCYC6-OO               C   7H  13O   2     G    300.00   4000.00 1386.00      1
 .252650839E+02 .325458915E-01-.113494502E-04 .178540172E-08-.104551384E-12    2
-.262255150E+05-.112686720E+03-.606776148E+01 .998265984E-01-.637962761E-04    3
 .191011484E-07-.207496071E-11-.148337709E+05 .575547331E+02                   4
MCYC6T-QOOH             C   7H  13O   2     G    300.00   4000.00 2055.00      1
 .234331685E+02 .347621964E-01-.124048044E-04 .199225952E-08-.118633947E-12    2
-.195868561E+05-.990888361E+02-.694095755E+01 .104651350E+00-.698281467E-04    3
 .219897276E-07-.260222584E-11-.958151058E+04 .634587763E+02                   4
MCYC6-OOQOOH            C   7H  13O   4     G    300.00   4000.00 1394.00      1
 .305321225E+02 .326136355E-01-.113442944E-04 .178165385E-08-.104214977E-12    2
-.403458401E+05-.135302325E+03-.434829022E+01 .112403701E+00-.796910207E-04    3
 .277878216E-07-.380650779E-11-.281870009E+05 .524217373E+02                   4
MCYC6T-OOQOOH           C   7H  13O   4     G    300.00   4000.00 1394.00      1
 .305321225E+02 .326136355E-01-.113442944E-04 .178165385E-08-.104214977E-12    2
-.403458401E+05-.135302325E+03-.434829022E+01 .112403701E+00-.796910207E-04    3
 .277878216E-07-.380650779E-11-.281870009E+05 .524217373E+02                   4
NC7H15                  C   7H  15          G    300.00   4000.00 1382.00      1
 .216371448E+02 .323324804E-01-.109273807E-04 .168357060E-08-.971774091E-13    2
-.105877217E+05-.852228493E+02-.379155767E-01 .756726570E-01-.407473634E-04    3
 .932678943E-08-.492360745E-12-.235605303E+04 .337321506E+02                   4
NC7H15-OO               C   7H  15O   2     G    300.00   4000.00 1393.00      1
 .272928290E+02 .327034748E-01-.112483701E-04 .175282538E-08-.101955579E-12    2
-.235449480E+05-.109307876E+03 .137396160E+01 .925294066E-01-.644403647E-04    3
 .235223293E-07-.356678305E-11-.144154775E+05 .302419431E+02                   4
NC7-QOOH                C   7H  15O   2     G    300.00   4000.00 1000.00      1
 .449365222E+02 .384325070E-02-.181753210E-06-.116055420E-10 .168632530E-14    2
-.301866739E+05-.207157897E+03 .169959950E+01 .943723540E-01-.755904260E-04    3
 .401131540E-07-.120065810E-10-.147076150E+05 .283145640E+02                   4
NC7-OOQOOH              C   7H  15O   4     G    300.00   4000.00 1395.00      1
 .269436049E+02 .351661203E-01-.120111248E-04 .186268617E-08-.107974911E-12    2
-.478858130E+05-.104588181E+03 .234060326E+01 .923428863E-01-.637138459E-04    3
 .236026902E-07-.368902757E-11-.392112217E+05 .278171493E+02                   4
!C6H4C2H                 C   8H   5          G    300.00   4000.00 1000.00      1 !polimi
! .286860656E+02-.138698600E-01 .227211900E-04-.998822700E-08 .140859000E-11    2
! .560473490E+05-.127502636E+03-.293242200E+01 .660436800E-01-.395005000E-04    3
!-.318303810E-08 .853003870E-11 .653240430E+05 .380586850E+02                   4
C6H4C2H C6H4-CCH  T10/13C  8.H  5.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.51356812E+01 1.95393656E-02-7.04783919E-06 1.14147499E-09-6.85061656E-14    2
 6.04891517E+04-5.42442195E+01-6.76311844E-01 5.42227756E-02-1.44506489E-05    3
-2.83755064E-08 1.79798680E-11 6.51966135E+04 2.93260540E+01 6.72297466E+04    4
!C6H5C2H2                C   8H   7          G    300.00   4000.00 1394.00      1 !Polimi
! .187667289E+02 .200619262E-01-.690883699E-05 .107799789E-08-.627759176E-13    2
! .376789029E+05-.760287256E+02-.272251268E+01 .709701368E-01-.527526320E-04    3
! .197369835E-07-.295890798E-11 .450007235E+05 .390143531E+02                   4
C6H5C2H2 n-styryl T12/07C  8.H  7.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.60668682E+01 2.35522834E-02-8.47352807E-06 1.36928204E-09-8.20829942E-14    2
 3.98109546E+04-6.01469382E+01 2.78678850E-01 4.12517677E-02 4.27417783E-05    3
-9.66212597E-08 4.47818574E-11 4.52024803E+04 2.70544015E+01 4.73269020E+04    4
!RXYLENE                 C   8H   9          G    300.00   4000.00 1000.00      1
! .808697123E+01 .442230490E-01-.196920930E-04 .391313300E-08-.286780230E-12    2
! .152828351E+05-.180507988E+02-.244083000E+01 .750206000E-01-.520941000E-04    3
! .184357000E-07-.267709000E-11 .180599500E+05 .358328500E+02                   4
RXYLENE           T 9/13C  8.H  9.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik  2-3C6H4CH2*
 1.56947853E+01 2.95619506E-02-1.06097584E-05 1.71214533E-09-1.02481459E-13    2
 1.41477221E+04-5.99627856E+01 5.72547012E-01 4.45565169E-02 4.13301302E-05    3
-9.20754733E-08 4.18729206E-11 1.95112053E+04 2.43021144E+01 2.18652673E+04    4
!C6H5CHCH3               C   8H   9          G    300.00   4000.00 1000.00      1 !EBenz old polimi
! .179749910E+02 .239625180E-01-.715492520E-05 .103757720E-08-.596944840E-13    2
! .194242850E+05-.693345570E+02-.526520200E+01 .889877600E-01-.754492360E-04    3
! .341497320E-07-.666954430E-11 .259605610E+05 .509400020E+02                   4
C6H5CHCH3 A1CHCH3 T 1/14C  8.H  9.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.52771567E+01 2.96305787E-02-1.06968599E-05 1.72910274E-09-1.03530176E-13    2
 1.47917666E+04-5.54929193E+01 2.27328453E+00 3.30022851E-02 6.58045139E-05    3
-1.15196192E-07 4.99525562E-11 1.98294339E+04 1.91733305E+01 2.23513746E+04    4
C6H5C2H4 A1CH2CH2* 11/04C  8.H  9.   0.   0.G   200.000  6000.000 1000.        1 !Burcat kik. ER add this species in PAH1906
 1.61326962E+01 2.82904273E-02-1.01801876E-05 1.64176637E-09-9.81375329E-14    2
 2.08791061E+04-6.00115413E+01 7.33299107E-01 4.59053158E-02 3.78257231E-05    3
-9.12367411E-08 4.25589678E-11 2.61572945E+04 2.50411074E+01 2.85902549E+04    4
C18H14 C9H7C9H7         H  14C  18          G   100.000  5000.000  990.27      1  !Kik add from Jin Hanfeng Combustion and Flame 206 (2019): 1-20.
 3.20125595E+01 5.89532847E-02-2.32102353E-05 4.57752278E-09-3.44228657E-13    2
 2.23209936E+04-1.51408560E+02-1.99662811E+00 8.71499057E-02 9.94525782E-05    3
-1.89332690E-07 7.67158406E-11 3.44098058E+04 3.93622783E+01                   4
RUME7                   C   8H  13O   2     G    300.00   4000.00 1376.00      1
 .270534591E+02 .305004468E-01-.106520501E-04 .167796515E-08-.983020287E-13    2
-.363346010E+05-.107800076E+03 .366021323E+01 .765652941E-01-.421034444E-04    3
 .990005395E-08-.618141131E-12-.272971814E+05 .209764369E+02                   4
RME7                    C   8H  15O   2     G    300.00   4000.00 1382.00      1
 .283088733E+02 .346001847E-01-.117889297E-04 .182346779E-08-.105527368E-12    2
-.507031223E+05-.115791454E+03 .312712425E+01 .886538094E-01-.550709022E-04    3
 .172495936E-07-.218153163E-11-.414147165E+05 .212562509E+02                   4
IC8H17                  C   8H  17          G    300.00   4000.00 1000.00      1
 .210071027E+02 .400670210E-01-.122220840E-04 .179139180E-08-.103364050E-12    2
-.156827594E+05-.841376688E+02-.142527150E+01 .952433870E-01-.515412500E-04    3
 .269038680E-08 .557281520E-11-.909216410E+04 .335841900E+02                   4
IC8-QOOH                C   8H  17O   2     G    300.00   4000.00 1400.00      1
 .323288504E+02 .354286616E-01-.121434812E-04 .188811322E-08-.109661472E-12    2
-.319868602E+05-.136609837E+03-.150530420E+01 .118500203E+00-.910186246E-04    3
 .362481173E-07-.587667874E-11-.206807572E+05 .436006519E+02                   4
IC8H17-OO               C   8H  17O   2     G    300.00   4000.00 1397.00      1
 .307492955E+02 .368544999E-01-.126522533E-04 .196915974E-08-.114442369E-12    2
-.380116818E+05-.129042218E+03-.126574300E+01 .113828908E+00-.844050615E-04    3
 .328104935E-07-.525271208E-11-.270886887E+05 .421608430E+02                   4
IC8T-QOOH               C   8H  17O   2     G    300.00   4000.00 1400.00      1
 .323288504E+02 .354286616E-01-.121434812E-04 .188811322E-08-.109661472E-12    2
-.319868602E+05-.136609837E+03-.150530420E+01 .118500203E+00-.910186246E-04    3
 .362481173E-07-.587667874E-11-.206807572E+05 .436006519E+02                   4
IC8-OOQOOH              C   8H  17O   4     G    300.00   4000.00 1398.00      1
 .362956073E+02 .372755603E-01-.128091685E-04 .199516372E-08-.116026947E-12    2
-.507708950E+05-.153592254E+03 .134208862E+01 .119507370E+00-.864939904E-04    3
 .319097725E-07-.475802942E-11-.387629197E+05 .338018650E+02                   4
!INDENYL                 C   9H   7          G    300.00   4000.00 1389.00      1 !polimi
! .210619876E+02 .219045968E-01-.772700080E-05 .122481766E-08-.721012249E-13    2
! .270100509E+05-.947705468E+02-.627808779E+01 .881610767E-01-.698280991E-04    3
! .280009421E-07-.454051640E-11 .362473103E+05 .511874555E+02                   4
!INDENYL           T 9/96C  9.H  7.   0.   0.G   200.000  6000.000  1000.       1 !Burcat kik 1-indenyl
! 1.85549761E+01 2.50350502E-02-9.14573755E-06 1.49348099E-09-9.01328268E-14    2
! 2.57211482E+04-7.63004782E+01-2.66986010E+00 6.21770959E-02 1.50674040E-05    3
!-7.96461960E-08 4.09191931E-11 3.23869684E+04 3.78611069E+01 3.43495696E+04    4
INDENYL           --G3B3H   7C   9          G     300.0    4000.0  1000.0    0 1  !AN 2100 from Jin at al 2019   10.1016/j.combustflame.2019.04.040
   1.40925252E1  3.36504564E-2  -1.5073094E-5  3.15831565E-9-2.52938691E-13    2
   2.65973353E4  -5.32839911E1  -1.19141936E1  1.27380531E-1   -1.554866E-4    3
  1.06821981E-7-3.12264529E-11   3.28223057E4   7.60295607E1                   4
RC9H11                  C   9H  11          G    300.00   4000.00 1385.00      1
 .227307929E+02 .291439937E-01-.101635526E-04 .159859987E-08-.935933623E-13    2
 .481056390E+04-.975266902E+02-.180604559E+01 .826070356E-01-.539943357E-04    3
 .177716542E-07-.237645289E-11 .137819561E+05 .357292291E+02                   4
!C10H7                   C  10H   7          G    300.00   4000.00 1000.00      1 !polimi
! .146529084E+02 .356159360E-01-.121796480E-04 .138747960E-08 .000000000E+00    2
! .405898415E+05-.575649187E+02-.631700500E+01 .913910790E-01-.608201990E-04    3
! .152228010E-07 .000000000E+00 .464268700E+05 .512234700E+02                   4
C10H7 Naphtyl rad T 7/98C  10H   7    0    0G   200.000  6000.000 1000.        1 !Burcat kik
 1.83535073E+01 2.77474314E-02-1.00885968E-05 1.64229575E-09-9.89002001E-14    2
 3.89261241E+04-7.48978150E+01-1.89559772E+00 5.83077290E-02 2.79388931E-05    3
-9.14375172E-08 4.46422302E-11 4.55409775E+04 3.52453263E+01 4.76546183E+04    4
!C10H7O                  C  10H   7O   1     G    300.00   4000.00 1387.00      1 !polimi
! .252263199E+02 .234793777E-01-.827533154E-05 .131107385E-08-.771548491E-13    2
! .188945294E+04-.112699321E+03-.234081413E+01 .850055448E-01-.590412510E-04    3
! .195981954E-07-.248272174E-11 .116463286E+05 .362009562E+02                   4
C10H7O    Radical T 7/98C 10.H  7.O  1.   0.G   200.000  6000.000 1000.00      1 !Burcat kik
 2.10591364E+01 2.82563070E-02-1.03328686E-05 1.68867034E-09-1.01974767E-13    2
 4.09143507E+03-8.84963398E+01-1.15176448E+00 6.11354512E-02 3.20151083E-05    3
-9.94285290E-08 4.79990043E-11 1.14058756E+04 3.25584836E+01 1.38887800E+04    4
C10H6OH   Radical T 7/98C 10.H  7.O  1.   0.G   200.000  6000.000 1000.00      1 !AN 2100 as C10H7O to be checked 
 2.10591364E+01 2.82563070E-02-1.03328686E-05 1.68867034E-09-1.01974767E-13    2
 4.09143507E+03-8.84963398E+01-1.15176448E+00 6.11354512E-02 3.20151083E-05    3
-9.94285290E-08 4.79990043E-11 1.14058756E+04 3.25584836E+01 1.38887800E+04    4
RTETRALIN               C  10H  11          G    300.00   4000.00 1393.00      1
 .274897602E+02 .290231662E-01-.101643070E-04 .160474752E-08-.942455736E-13    2
 .498834588E+04-.134140516E+03-.103201226E+02 .112759920E+00-.777366610E-04    3
 .248527119E-07-.289510552E-11 .183518811E+05 .701782401E+02                   4
RTETRAOO                C  10H  11O   2     G    300.00   4000.00 1393.00      1
 .325696052E+02 .270322587E-01-.103226960E-04 .172977036E-08-.105947326E-12    2
-.797598133E+04-.153101057E+03-.133437809E+02 .139730780E+00-.110918062E-03    3
 .406822937E-07-.565600132E-11 .639529388E+04 .899902305E+02                   4
RODECA                  C  10H  17          G    300.00   4000.00 1393.00      1
 .266885367E+02 .438181872E-01-.149997894E-04 .233096426E-08-.135354849E-12    2
-.142864228E+05-.128706101E+03-.137726588E+02 .134621624E+00-.905467076E-04    3
 .298633466E-07-.381482514E-11-.121358784E+02 .896659972E+02                   4
RDECALIN                C  10H  17          G    300.00   4000.00 1393.00      1
 .266885367E+02 .438181872E-01-.149997894E-04 .233096426E-08-.135354849E-12    2
-.142864228E+05-.128706101E+03-.137726588E+02 .134621624E+00-.905467076E-04    3
 .298633466E-07-.381482514E-11-.121358784E+02 .896659972E+02                   4
RDECOO                  C  10H  17O   2     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
QDECOOH                 C  10H  17O   2     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
ZDECA                   C  10H  17O   4     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
NC10H19                 C  10H  19          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC10H21                 C  10H  21          G    300.00   4000.00 1385.00      1
 .314447580E+02 .452778532E-01-.153145696E-04 .236072411E-08-.136311835E-12    2
-.229702700E+05-.131435127E+03-.930536886E+00 .113137924E+00-.664034118E-04    3
 .183220872E-07-.177128003E-11-.109890165E+05 .451328034E+02                   4
NC10-QOOH               C  10H  21O   2     G    300.00   4000.00 1392.00      1
 .364873664E+02 .456938220E-01-.154604572E-04 .238346695E-08-.137626430E-12    2
-.370093465E+05-.152798812E+03 .883511244E+00 .125360621E+00-.820308363E-04    3
 .270294818E-07-.354081617E-11-.243570772E+05 .395546233E+02                   4
NC10H21-OO              C  10H  21O   2     G    300.00   4000.00 1392.00      1
 .347424373E+02 .481682266E-01-.165183738E-04 .256870455E-08-.149189141E-12    2
-.416206773E+05-.145293449E+03 .109633829E+01 .123998092E+00-.822926235E-04    3
 .288935474E-07-.426829326E-11-.295195291E+05 .366210584E+02                   4
NC10-OOQOOH             C  10H  21O   4     G    300.00   4000.00 1393.00      1
 .419701067E+02 .470326141E-01-.162065055E-04 .252885796E-08-.147242779E-12    2
-.568721943E+05-.179987435E+03 .270340236E+01 .134161981E+00-.884509572E-04    3
 .291143638E-07-.380678318E-11-.428023111E+05 .324857210E+02                   4
!C10H7CH2                C  11H   9          G    300.00   4000.00 1389.00      1 !polimi
! .266596927E+02 .269903845E-01-.949827903E-05 .150313533E-08-.883831941E-13    2
! .210179470E+05-.122975754E+03-.551514480E+01 .106245066E+00-.857510752E-04    3
! .355122444E-07-.598055713E-11 .318146452E+05 .484291679E+02                   4
C10H7CH2          T 7/98C  11H   9    0    0G   200.000  6000.000 1000.        1 !Burcat kik 1-C10H7-CH2*
 2.18977539E+01 3.26102636E-02-1.18401218E-05 1.92574628E-09-1.15903442E-13    2
 2.24571098E+04-9.41050741E+01-2.53234304E+00 7.32920338E-02 2.02974707E-05    3
-9.36547823E-08 4.70753594E-11 3.02906705E+04 3.79638513E+01 3.28097266E+04    4
!C10H6CH3                C  11H   9          G    300.00   4000.00 1387.00      1 !polimi
! .241866524E+02 .287085863E-01-.100040198E-04 .157283341E-08-.920615442E-13    2
! .317595121E+05-.107209439E+03-.148986180E+01 .837301572E-01-.531437515E-04    3
! .161159556E-07-.183550466E-11 .411521411E+05 .324161445E+02                   4
C10H6CH3          T11/13C 11.H  9.   0.   0.G   200.000  6000.000  1000.       1 !burcat kik 1-Naphthyl-3-Methyl Radical 1-C10H6*-3-CH3 
 2.06757697E+01 3.29978114E-02-1.19213860E-05 1.93272353E-09-1.16069177E-13    2
 3.42587802E+04-8.79526119E+01-2.07498418E+00 6.80090538E-02 2.63761043E-05    3
-9.53060559E-08 4.65647314E-11 4.17116175E+04 3.57867673E+01 4.41824233E+04    4
CH3C10H6O               C  11H   9O   1     G    300.00   4000.00 1386.00      1
 .281108749E+02 .281427040E-01-.986090177E-05 .155620703E-08-.913337710E-13    2
-.350666986E+04-.125748079E+03-.108570461E+01 .905308669E-01-.577474885E-04    3
 .167977934E-07-.168045736E-11 .709977655E+04 .329292729E+02                   4
O2C10H6CH3              C  11H   9O   2     G    200.00   3500.00 1000.00      1 !AN 2100
 1.35895989e+01 5.87348211e-02-3.12371840e-05 7.93473778e-09-7.75713505e-13    2
 1.23461692e+04-4.57265893e+01-1.41546285e+01 1.69711731e-01-1.97702548e-04    3
 1.18911647e-07-2.85199409e-11 1.78950146e+04 8.81232703e+01                   4
C10H7CH2OOH             C  11H  10O   2     G    200.00   3500.00 1000.00      1 !AN 2100
 9.59357138e+00 7.25131650e-02-4.02299436e-05 1.04419276e-08-1.03126751e-12    2
-1.67373550e+03-1.93308190e+01-1.20905038e+01 1.59249466e-01-1.70334395e-04    3
 9.71782283e-08-2.27153427e-11 2.66307953e+03 8.52823091e+01                   4
OC10H6CH2               C  11H   8O   1     G    200.00   3500.00 1190.00      1 !AN 2100
 1.61060825e+01 4.46337369e-02-2.08038137e-05 4.64415651e-09-4.06679510e-13    2
 5.08234293e+03-6.36614858e+01-1.01446499e+01 1.32871493e-01-1.32027876e-04    3
 6.69545554e-08-1.34970994e-11 1.13300172e+04 6.75495253e+01                   4
C10H7CH2O               C  11H   9O   1     G    200.00   3500.00 1000.00      1 !AN 2100
 6.19208112e+00 6.85969273e-02-3.75702665e-05 9.69725993e-09-9.55827851e-13    2
 1.63598794e+04-4.97892094e+00-1.25750275e+01 1.43665362e-01-1.50172918e-04    3
 8.47656942e-08-1.97229364e-11 2.01133012e+04 8.55615295e+01                   4
C10H7CH2O2              C  11H   9O   2     G    200.00   3500.00 1000.00      1 !AN 2100
 1.10033962e+01 6.55567635e-02-3.57758606e-05 9.18803899e-09-9.01110330e-13    2
 1.54881793e+04-2.80172408e+01-1.29736639e+01 1.61465004e-01-1.79638221e-04    3
 1.05096279e-07-2.48781704e-11 2.02835913e+04 8.76582139e+01                   4
RUME10                  C  11H  19O   2     G    300.00   4000.00 1400.00      1
 .333201898E+02 .479399831E-01-.157699228E-04 .238393079E-08-.135735725E-12    2
-.400970534E+05-.137405141E+03 .142231026E+01 .127120401E+00-.922642215E-04    3
 .364453822E-07-.599028369E-11-.294852312E+05 .322500169E+02                   4
RMDX                    C  11H  21O   2     G    300.00   4000.00 1376.00      1
 .385051195E+02 .464902832E-01-.162008540E-04 .254969816E-08-.149299808E-12    2
-.649901621E+05-.166525707E+03 .345128941E+01 .114960511E+00-.621890037E-04    3
 .140937438E-07-.752795690E-12-.513892174E+05 .266431624E+02                   4
QMDOOH                  C  11H  21O   4     G    300.00   4000.00 1378.00      1
 .463512360E+02 .442905004E-01-.156791241E-04 .249437540E-08-.147109263E-12    2
-.802179278E+05-.202701285E+03 .505901193E+01 .130586874E+00-.811966955E-04    3
 .236808295E-07-.254638441E-11-.648189073E+05 .227472201E+02                   4
RMDOOX                  C  11H  21O   4     G    300.00   4000.00 1384.00      1
 .426675367E+02 .481355870E-01-.164385340E-04 .254942818E-08-.147838407E-12    2
-.850035553E+05-.184014175E+03 .443641793E+01 .133210481E+00-.883606205E-04    3
 .302231077E-07-.426647212E-11-.712160785E+05 .229630078E+02                   4
ZMDOOH                  C  11H  21O   6     G    300.00   4000.00 1384.00      1
 .493171232E+02 .461887725E-01-.155948619E-04 .242596048E-08-.141314237E-12    2
-.997314376E+05-.213131636E+03 .613115269E+01 .145831804E+00-.103807590E-03    3
 .382530920E-07-.579145154E-11-.845666547E+05 .193222210E+02                   4
!C12H7                   C  12H   7          G    300.00   4000.00 1000.00      1 !polimi
! .119534365E+02 .523860720E-01-.276952580E-04 .698583900E-08-.684938540E-12    2
! .531995141E+05-.403925438E+02-.733802700E+01 .111965800E+00-.932829430E-04    3
! .358663430E-07-.426602200E-11 .580597660E+05 .573507160E+02                   4
C12H7 AcenaphtynylT01/08C 12.H  7.   0.   0.G   200.000  6000.000  1000.00     1 !Burcat kik
 2.16586138E+01 3.04696316E-02-1.11497201E-05 1.82316781E-09-1.10144488E-13    2
 5.28451416E+04-9.73300058E+01-2.23704309E+00 6.20074173E-02 4.69635631E-05    3
-1.20874263E-07 5.68318739E-11 6.08867652E+04 3.38045560E+01 6.31787081E+04    4
!C12H9                       C  12H   9          G    300.00   4000.00 1000.00      1 !polimi
! .214890352E+02 .375797860E-01-.121080230E-04 .129882780E-08 .000000000E+00    2
! .415521488E+05-.916763235E+02-.783196500E+01 .114327200E+00-.776398370E-04    3
! .194042280E-07 .000000000E+00 .498170300E+05 .608493300E+02                   4
C12H9                   C  12H   9          G    300.00   6000.00 1000.00      1 !Burcat kik P2-
 2.25692222E+01 3.45619984E-02-1.27020877E-05 2.08111819E-09-1.25849407E-13    2
 4.05907457E+04-9.57787051E+01 4.07668089E-01 5.42794698E-02 7.12515775E-05    3
-1.44404112E-07 6.48497982E-11 4.85351870E+04 2.81980814E+01 5.14438013E+04    4
NC12H25                 C  12H  25          G    300.00   4000.00 1387.00      1
 .379559371E+02 .541231481E-01-.184408520E-04 .285618139E-08-.165452331E-12    2
-.312698454E+05-.166157365E+03-.117025753E+01 .136564242E+00-.813840519E-04    3
 .231564976E-07-.240764498E-11-.167979250E+05 .471339366E+02                   4
NC12-QOOH               C  12H  25O   2     G    300.00   4000.00 1392.00      1
 .427882927E+02 .547351985E-01-.185693137E-04 .286771608E-08-.165782124E-12    2
-.451897912E+05-.183774591E+03 .457142729E+00 .149660990E+00-.984019129E-04    3
 .327982507E-07-.438634589E-11-.301386488E+05 .448987214E+02                   4
NC12H25-OO              C  12H  25O   2     G    300.00   4000.00 1392.00      1
 .410672882E+02 .571682582E-01-.196096581E-04 .304996352E-08-.177163659E-12    2
-.498119415E+05-.176403781E+03 .761653139E+00 .147870053E+00-.980093227E-04    3
 .342486611E-07-.502171364E-11-.353144020E+05 .415448990E+02                   4
NC12-OOQOOH             C  12H  25O   4     G    300.00   4000.00 1393.00      1
 .478223133E+02 .563342752E-01-.193784199E-04 .302016363E-08-.175696376E-12    2
-.648031378E+05-.208209874E+03 .250560092E+01 .157994999E+00-.105503812E-03    3
 .358709948E-07-.494871123E-11-.486270464E+05 .366890378E+02                   4
!C14H9                   C  14H   9          G    300.00   4000.00 1000.00      1 !polimi
! .255171870E+02 .393727940E-01-.123155080E-04 .127852800E-08 .000000000E+00    2
! .431324738E+05-.115618425E+03-.909474100E+01 .131333800E+00-.924017290E-04    3
! .240156710E-07 .000000000E+00 .527750200E+05 .639753600E+02                   4
C14H9 4-Phenantr  T11/07C 14.H  9.   0.   0.G   298.150  5000.000  1000.00     1 !Burcat kik assume 4-Phenanthryl rad as it is active site to from pyrene
 2.68173412E+01 3.76935761E-02-1.45586251E-05 2.58486800E-09-1.73198001E-13    2
 4.14405846E+04-1.21547559E+02-1.08929968E+01 1.41537035E-01-1.14205532E-04    3
 3.57710437E-08 0.00000000E+00 5.21136455E+04 7.37137024E+01 5.42184687E+04    4
C16H9                   C  16H   9          G    300.00   4000.00 1000.00      1
 .161628784E+02 .696969850E-01-.371786410E-04 .946306230E-08-.935417110E-12    2
 .461067047E+05-.652717249E+02-.114972670E+02 .151166960E+00-.116351410E-03    3
 .317097570E-07 .218082760E-11 .532378630E+05 .757195740E+02                   4
C18H9                   C  18H   9          G    300.00   3500.00 1240.00      1 !test C18H9=C16H9+(C16H9-C14H9)
 7.28131520E+00 9.79858540E-02-5.71014164E-05 1.55232196E-08-1.60913985E-12    2
 5.01527171E+04-1.86201194E+01-1.50799037E+01 1.82129796E-01-1.71943851E-04    3
 8.35734254E-08-1.64715049E-11 5.46706402E+04 9.01438864E+01                   4
!C18H9                   C  18H   9          G    300.00   4000.00 1000.00      1     !KS 1800
! 6.80856980E+00	1.00021180E-01-6.20417740E-05	1.76475970E-08-1.8708342E-12     2
! 1.35345880E+05-2.46161870E+02-1.38997900E+01	1.71000120E-01-1.4030109E-04     3
! 3.94038430E-08	4.36165520E-12 5.37007060E+04	8.74637880E+01                   4
IC16H33                 C  16H  33          G    300.00   4000.00 1398.00      1
 .560389730E+02 .668182464E-01-.225681513E-04 .347608102E-08-.200620637E-12    2
-.583645424E+05-.270643351E+03-.953227198E+01 .224283987E+00-.166371012E-03    3
 .627848165E-07-.951119300E-11-.362947496E+05 .795385858E+02                   4
NC16H33                 C  16H  33          G    300.00   4000.00 1387.00      1
 .510324990E+02 .711045684E-01-.240491592E-04 .370710805E-08-.214054039E-12    2
-.477151440E+05-.228063103E+03-.243005348E+01 .186692969E+00-.115724867E-03    3
 .350879669E-07-.405848895E-11-.282942913E+05 .622394761E+02                   4
IC16H33-OO              C  16H  33O   2     G    300.00   4000.00 1397.00      1
 .600009189E+02 .697612153E-01-.240119992E-04 .374399505E-08-.217877031E-12    2
-.771125672E+05-.288496873E+03-.807177622E+01 .238256241E+00-.186291159E-03    3
 .758296536E-07-.125956694E-10-.544214916E+05 .737310481E+02                   4
NC16-QOOH               C  16H  33O   2     G    300.00   4000.00 1394.00      1
 .557196631E+02 .758805933E-01-.260092776E-04 .404350192E-08-.234807139E-12    2
-.852319237E+05-.250905152E+03-.858601178E+00 .204663464E+00-.138309577E-03    3
 .488963438E-07-.717831502E-11-.651200924E+05 .543621098E+02                   4
IC16-QOOH               C  16H  33O   2     G    300.00   4000.00 1399.00      1
 .615798034E+02 .683372119E-01-.235040286E-04 .366308625E-08-.213104512E-12    2
-.710887760E+05-.294961987E+03-.836284759E+01 .243137667E+00-.193204766E-03    3
 .794478202E-07-.132585716E-10-.480052296E+05 .765156723E+02                   4
NC16H33-OO              C  16H  33O   2     G    300.00   4000.00 1392.00      1
 .537254976E+02 .751675700E-01-.257930312E-04 .401271756E-08-.233130903E-12    2
-.661992854E+05-.238675214E+03 .121036107E+00 .195526928E+00-.129332034E-03    3
 .448994551E-07-.651714304E-11-.469097176E+05 .512502917E+02                   4
IC16T-QOOH              C  16H  33O   2     G    300.00   4000.00 1397.00      1
 .619590914E+02 .670805941E-01-.228781110E-04 .354645272E-08-.205581639E-12    2
-.737750910E+05-.297686975E+03-.828638110E+01 .240615134E+00-.188046280E-03    3
 .753924180E-07-.122092604E-10-.505105835E+05 .759168895E+02                   4
IC16T-OOQOOH            C  16H  33O   4     G    300.00   4000.00 1396.00      1
 .664600695E+02 .692200495E-01-.239811044E-04 .375550159E-08-.219211037E-12    2
-.927495777E+05-.318609160E+03-.734744585E+01 .256652224E+00-.210530384E-03    3
 .896944245E-07-.155165690E-10-.685533247E+05 .725686554E+02                   4
NC16-OOQOOH             C  16H  33O   4     G    300.00   4000.00 1393.00      1
 .605564321E+02 .743085731E-01-.255622121E-04 .398394439E-08-.231762903E-12    2
-.812450313E+05-.270973587E+03 .185761468E+01 .205470409E+00-.136236709E-03    3
 .460471713E-07-.632675050E-11-.602164277E+05 .464682670E+02                   4
IC16-OOQOOH             C  16H  33O   4     G    300.00   4000.00 1395.00      1
 .657312368E+02 .698159219E-01-.241818212E-04 .378635278E-08-.220988765E-12    2
-.891725518E+05-.313140345E+03-.709314164E+01 .252307521E+00-.202956898E-03    3
 .848048060E-07-.144255682E-10-.650715559E+05 .736645741E+02                   4
RUME16                  C  17H  31O   2     G    300.00   4000.00 1836.00      1
 .492312959E+02 .809629787E-01-.290414743E-04 .466984560E-08-.277987170E-12    2
-.712766099E+05-.212350222E+03 .581847898E+00 .197335153E+00-.132222747E-03    3
 .454132116E-07-.638160297E-11-.555076491E+05 .468001664E+02                   4
RMPAX                   C  17H  33O   2     G    300.00   4000.00 1000.00      1
 .347969412E+02 .108174887E+00-.436560662E-04 .805036686E-08-.557001848E-12    2
-.833532968E+05-.136711346E+03 .118429649E+02 .108281798E+00 .937470576E-04    3
-.175260710E-06 .681980157E-10-.741770519E+05-.304443036E+01                   4
RMPAOOX                 C  17H  33O   4     G    300.00   4000.00 1384.00      1
 .426675367E+02 .481355870E-01-.164385340E-04 .254942818E-08-.147838407E-12    2
-.850035553E+05-.184014175E+03 .443641793E+01 .133210481E+00-.883606205E-04    3
 .302231077E-07-.426647212E-11-.712160785E+05 .229630078E+02                   4
QMPAOOH                 C  17H  33O   4     G    300.00   4000.00 1378.00      1
 .463512360E+02 .442905004E-01-.156791241E-04 .249437540E-08-.147109263E-12    2
-.802179278E+05-.202701285E+03 .505901193E+01 .130586874E+00-.811966955E-04    3
 .236808295E-07-.254638441E-11-.648189073E+05 .227472201E+02                   4
ZMPAOOH                 C  17H  33O   6     G    300.00   4000.00 1384.00      1
 .493171232E+02 .461887725E-01-.155948619E-04 .242596048E-08-.141314237E-12    2
-.997314376E+05-.213131636E+03 .613115269E+01 .145831804E+00-.103807590E-03    3
 .382530920E-07-.579145154E-11-.845666547E+05 .193222210E+02                   4
RMLIN1X                 C  19H  31O   2     G    300.00   4000.00 1830.00      1
 .515951901E+02 .848982968E-01-.306132424E-04 .493978264E-08-.294767670E-12    2
-.437090861E+05-.222319284E+03-.124182769E+01 .210470141E+00-.141012967E-03    3
 .480938977E-07-.668889816E-11-.265018940E+05 .594297783E+02                   4
RMLIN1A                 C  19H  31O   2     G    300.00   4000.00 1830.00      1
 .515951901E+02 .848982968E-01-.306132424E-04 .493978264E-08-.294767670E-12    2
-.437090861E+05-.222319284E+03-.124182769E+01 .210470141E+00-.141012967E-03    3
 .480938977E-07-.668889816E-11-.265018940E+05 .594297783E+02                   4
RMLIN1OOX               C  19H  31O   4     G    300.00   4000.00 1854.00      1
 .566771062E+02 .848718923E-01-.306165992E-04 .494186779E-08-.294961213E-12    2
-.712260452E+05-.243221478E+03-.182318626E+01 .229267759E+00-.163619600E-03    3
 .597071790E-07-.884702825E-11-.526983896E+05 .668009912E+02                   4
QMLIN1OOX               C  19H  31O   4     G    300.00   4000.00 1859.00      1
 .597198037E+02 .825172318E-01-.298594827E-04 .482987333E-08-.288709215E-12    2
-.679692648E+05-.260058551E+03-.300959205E+01 .239625356E+00-.176824958E-03    3
 .662378545E-07-.999748235E-11-.483423909E+05 .715224170E+02                   4
ZMLIN1OOX               C  19H  31O   6     G    300.00   4000.00 1844.00      1
 .633953698E+02 .840133680E-01-.304696355E-04 .493592631E-08-.295352525E-12    2
-.861431583E+05-.275575442E+03 .377427203E+00 .239045319E+00-.172299424E-03    3
 .627369839E-07-.920510825E-11-.661691485E+05 .585014961E+02                   4
RMLINX                  C  19H  33O   2     G    300.00   4000.00 1386.00      1
 .611078575E+02 .762751735E-01-.262266430E-04 .408707626E-08-.237771674E-12    2
-.683962704E+05-.275956500E+03-.144781566E+01 .215019809E+00-.142192171E-03    3
 .476963895E-07-.649336150E-11-.458716461E+05 .627347784E+02                   4
RMLINA                  C  19H  33O   2     G    300.00   4000.00 1386.00      1
 .611078575E+02 .762751735E-01-.262266430E-04 .408707626E-08-.237771674E-12    2
-.683962704E+05-.275956500E+03-.144781566E+01 .215019809E+00-.142192171E-03    3
 .476963895E-07-.649336150E-11-.458716461E+05 .627347784E+02                   4
RMLIN1OH                C  19H  33O   3     G    300.00   4000.00 1000.00      1
 .109866520E+03 .423976550E-02-.805195410E-07-.170406780E-10 .168247750E-14    2
-.106680810E+06-.543129330E+03 .690969590E+00 .209334020E+00-.125946550E-03    3
 .409375960E-07-.109953440E-10-.661363050E+05 .579650690E+02                   4
RMLINOOX                C  19H  33O   4     G    300.00   4000.00 1840.00      1
 .561396497E+02 .898573320E-01-.323076347E-04 .520295879E-08-.310043109E-12    2
-.835647272E+05-.240835194E+03 .146002415E+01 .221120424E+00-.149309126E-03    3
 .517229930E-07-.733489301E-11-.658774535E+05 .502873652E+02                   4
QMLINOOX                C  19H  33O   4     G    300.00   4000.00 1830.00      1
 .592334771E+02 .871071695E-01-.313329462E-04 .504827960E-08-.300945381E-12    2
-.780101129E+05-.256778117E+03-.383425349E+00 .231626065E+00-.160960610E-03    3
 .566395921E-07-.805109149E-11-.589322117E+05 .599912602E+02                   4
RMLIN1OHOO              C  19H  33O   5     G    300.00   4000.00 1000.00      1
 .251712040E+02 .137856480E+00-.512202200E-04 .870306320E-08-.560550030E-12    2
-.886761250E+05-.568400270E+02-.493498520E+01 .253526120E+00-.181310740E-03    3
 .532790980E-07-.715418010E-12-.841542810E+05 .856818080E+02                   4
ZMLINOOX                C  19H  33O   6     G    300.00   4000.00 1183.00      1
 .601829822E+02 .877246704E-01-.308673874E-04 .490011538E-08-.289106438E-12    2
-.959756017E+05-.274111539E+03 .888177201E+00 .245491279E+00-.188867182E-03    3
 .756398491E-07-.122061299E-10-.781464330E+05 .361650421E+02                   4
RMEOLEA                 C  19H  35O   2     G    300.00   4000.00 1386.00      1
 .617968812E+02 .797287018E-01-.272798012E-04 .423721781E-08-.245941529E-12    2
-.826622063E+05-.278715034E+03-.296860913E-01 .215538273E+00-.139084893E-03    3
 .453526106E-07-.596335185E-11-.602711250E+05 .564905254E+02                   4
RMEOLES                 C  19H  35O   2     G    300.00   4000.00 1386.00      1
 .617968812E+02 .797287018E-01-.272798012E-04 .423721781E-08-.245941529E-12    2
-.826622063E+05-.278715034E+03-.296860913E-01 .215538273E+00-.139084893E-03    3
 .453526106E-07-.596335185E-11-.602711250E+05 .564905254E+02                   4
RMEOLEOOX               C  19H  35O   4     G    300.00   4000.00 1799.00      1
 .565118676E+02 .949710722E-01-.342666750E-04 .553134168E-08-.330143553E-12    2
-.121723087E+06-.240377715E+03 .312228984E+01 .215930145E+00-.133878272E-03    3
 .413627115E-07-.514696341E-11-.103763030E+06 .464356398E+02                   4
QMEOLEOOH               C  19H  35O   4     G    300.00   4000.00 1825.00      1
 .578903822E+02 .960618008E-01-.345783142E-04 .557312937E-08-.332293982E-12    2
-.145787244E+06-.248797880E+03-.121085721E+01 .236084007E+00-.157011163E-03    3
 .530523572E-07-.729693062E-11-.126516243E+06 .664772594E+02                   4
ZMEOLEOOX               C  19H  35O   6     G    300.00   4000.00 1175.00      1
 .558298346E+02 .101939581E+00-.350749088E-04 .548251413E-08-.319925836E-12    2
-.108843753E+06-.228788516E+03 .196924109E+01 .244903891E+00-.177892306E-03    3
 .692918136E-07-.110530115E-10-.926192007E+05 .531689573E+02                   4
RSTEAX                  C  19H  37O   2     G    300.00   4000.00 1000.00      1
 .410838828E+02 .116388491E+00-.460844475E-04 .839784976E-08-.576703150E-12    2
-.912925804E+05-.167019971E+03 .115570681E+02 .131479341E+00 .799583356E-04    3
-.171755777E-06 .679701047E-10-.799964069E+05 .174630364E+01                   4
RMEOLEOH                C  19H  37O   3     G    300.00   4000.00 1000.00      1
 .113871410E+03 .775875800E-02-.452147480E-06 .136135370E-10-.133024960E-16    2
-.136912560E+06-.564887510E+03 .250303720E+01 .215053450E+00-.121530550E-03    3
 .330490980E-07-.788034390E-11-.955148750E+05 .486207620E+02                   4
QMSTEAOOH               C  19H  37O   4     G    300.00   3500.00 1230.00      1
-1.30612112e+02 6.00365407e-01-4.85197507e-04 1.58690694e-07-1.80918278e-11    2
 1.24045712e+04 7.12083733e+02 2.15554520e+01 1.05511541e-01 1.18282818e-04    3
-1.68398913e-07 4.83897995e-11-2.50286495e+04-5.35376428e+01                   4
RMSTEAOOX               C  19H  37O   4     G    300.00   3500.00 1250.00      1
-1.20700825e+02 5.67736647e-01-4.52750605e-04 1.47317719e-07-1.67528750e-11    2
 1.02039730e+04 6.60024010e+02 1.91170969e+01 1.20319296e-01 8.41502164e-05    3
-1.39029386e-07 4.05165459e-11-2.47505076e+04-4.57161098e+01                   4
RMEOLEOHOO              C  19H  37O   5     G    300.00   4000.00 1000.00      1
 .133736930E+02 .167858470E+00-.644862230E-04 .112143850E-07-.733979720E-12    2
-.112646060E+06 .973074340E+01-.366680260E+01 .261956100E+00-.180087150E-03    3
 .445610300E-07 .429013550E-11-.113462220E+06 .787735670E+02                   4
ZMSTEAOOH               C  19H  37O   6     G    300.00   3500.00 1250.00      1
-6.22995292e+01 3.41575945e-01-2.69706994e-04 8.71969173e-08-9.87435445e-12    2
 1.57160052e+04 3.57020399e+02 1.61954271e+01 9.03920846e-02 3.17136383e-05    3
-7.35607532e-08 2.22771796e-11-3.90773390e+03-3.91880337e+01                   4
!C10H8                   C  10H   8          G    300.00   4000.00 1401.00      1 !polimi
! .234023214E+02 .242434427E-01-.836282016E-05 .130620111E-08-.761153748E-13    2
! .651941329E+04-.107433208E+03-.883645988E+01 .109300567E+00-.955200914E-04    3
! .421647669E-07-.739851710E-11 .166533366E+05 .621064766E+02                   4
C10H8 Naphthalene T 7/98C  10H   8    0    0G   200.000  6000.000 1000.        1 !Burcat kik
 1.86129884E+01 3.04494175E-02-1.11224825E-05 1.81615474E-09-1.09601281E-13    2
 8.91578988E+03-8.00230396E+01-1.04919475E+00 4.62970781E-02 7.07591636E-05    3
-1.38408111E-07 6.20475407E-11 1.59848987E+04 3.02121626E+01 1.81107678E+04    4
NC3H7O2                 C   3H   7O   2     G    300.00   4000.00 1388.00      1
 .127230991E+02 .167336808E-01-.575943184E-05 .897769493E-09-.522275065E-13    2
-.108816595E+05-.381965321E+02 .156301709E+01 .426192697E-01-.296615075E-04    3
 .114187326E-07-.189894471E-11-.688086375E+04 .219842933E+02                   4
IC3H7O2                 C   3H   7O   2     G    300.00   4000.00 1392.00      1
 .132610651E+02 .162501084E-01-.558631798E-05 .870057473E-09-.505849469E-13    2
-.131937089E+05-.421023499E+02 .103495454E+01 .469942369E-01-.366525520E-04    3
 .157084173E-07-.281956117E-11-.906344820E+04 .229566921E+02                   4
NC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1374.00      1
 .146139980E+02 .143723015E-01-.488635144E-05 .756519620E-09-.438364992E-13    2
-.646101457E+04-.457478245E+02 .191005011E+01 .411666833E-01-.251630217E-04    3
 .711856873E-08-.698838732E-12-.179305093E+04 .234514457E+02                   4
IC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1399.00      1
 .155030898E+02 .139802008E-01-.481811216E-05 .751835399E-09-.437743118E-13    2
-.741643030E+04-.523911482E+02-.184042862E+00 .564670638E-01-.501611253E-04    3
 .230526863E-07-.423866481E-11-.252333896E+04 .298354826E+02                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1388.00      1
 .185146106E+02 .164157074E-01-.573085844E-05 .901975314E-09-.528299084E-13    2
-.231819444E+05-.618247164E+02 .254387733E+01 .570847379E-01-.472164204E-04    3
 .208289492E-07-.378162942E-11-.178600410E+05 .229447574E+02                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1391.00      1
 .191234208E+02 .158457151E-01-.552231946E-05 .868162288E-09-.508094203E-13    2
-.255253957E+05-.661419362E+02 .175906535E+01 .624712381E-01-.554930416E-04    3
 .257973727E-07-.483190839E-11-.200009572E+05 .251348546E+02                   4
CHOCH2CHO               C   3H   4O   2     G    300.00   4000.00 1000.00      1
 .104962923E+02 .120559957E-01-.434149310E-05 .699425892E-09-.418003976E-13    2
-.437332461E+05-.275425657E+02 .124227207E+01 .300698605E-01-.148206586E-05    3
-.242738150E-07 .133121686E-10-.408667843E+05 .219242842E+02                   4
C3H6O                   C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .801491079E+01 .173919953E-01-.626027968E-05 .101188256E-08-.606239111E-13    2
-.151980838E+05-.188279964E+02 .342806676E+01 .625176642E-02 .613196311E-04    3
-.860387185E-07 .351371393E-10-.128446646E+05 .104244994E+02                   4
NC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1000.00      1
 .852377408E+01 .210371210E-01-.748398370E-05 .119958663E-08-.714873013E-13    2
-.350702414E+05-.177857176E+02 .541877541E+01-.575566129E-03 .851215375E-04    3
-.111060442E-06 .443007063E-10-.328368377E+05 .529974117E+01                   4
IC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1000.00      1
 .964183701E+01 .200230715E-01-.711967189E-05 .114138950E-08-.679935249E-13    2
-.374835623E+05-.256288343E+02 .430755345E+01 .102582798E-01 .619565411E-04    3
-.902973802E-07 .373936384E-10-.349249212E+05 .755995822E+01                   4
C3H7OOH                 C   3H   8O   2     G    300.00   4000.00 1000.00      1
 .104115631E+02 .213763889E-01-.755819870E-05 .120207180E-08-.711798090E-13    2
-.268935445E+05-.235428789E+02 .708977756E+01-.486163264E-02 .103253531E-03    3
-.133200956E-06 .530799252E-10-.244194556E+05 .174859215E+01                   4
C3-OQOOH                C   3H   6O   3     G    300.00   4000.00 1391.00      1
 .170285271E+02 .130716784E-01-.459310856E-05 .726135156E-09-.426658337E-13    2
-.416334217E+05-.592513577E+02 .768933034E+00 .546905880E-01-.465072405E-04    3
 .203159585E-07-.358398999E-11-.363238861E+05 .268291637E+02                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   4000.00 1000.00      1
 .838041157E+01 .195206120E-01-.697374143E-05 .112144919E-08-.669467831E-13    2
-.848625211E+04-.189916219E+02 .421934640E+01 .738556641E-02 .602825529E-04    3
-.838680247E-07 .339623435E-10-.623491852E+04 .808139850E+01                   4
CH2OHCH2CHO             C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .118936666E+02 .144153203E-01-.477525443E-05 .726036430E-09-.415285995E-13    2
-.459271652E+05-.327285750E+02 .266613285E+01 .346302298E-01-.214380719E-04    3
 .690469334E-08-.916939105E-12-.425706030E+05 .173358364E+02                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   4000.00 1386.00      1
 .110500439E+02 .152562747E-01-.517257413E-05 .798146428E-09-.461030406E-13    2
-.142779432E+05-.312276095E+02 .149130595E+01 .376502110E-01-.258507542E-04    3
 .978662277E-08-.158835656E-11-.109017244E+05 .201908977E+02                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   4000.00 1388.00      1
 .110944203E+02 .153549108E-01-.523574640E-05 .810964124E-09-.469665855E-13    2
-.134769536E+05-.307070215E+02 .584672920E+00 .407370189E-01-.294865043E-04    3
 .116950656E-07-.196228356E-11-.984929391E+04 .255429190E+02                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   4000.00 1392.00      1
 .106573810E+02 .155684549E-01-.527663821E-05 .814099260E-09-.470228616E-13    2
-.112728087E+05-.272448749E+02 .975268381E+00 .369225253E-01-.232066980E-04    3
 .768472523E-08-.106762046E-11-.774554528E+04 .252661698E+02                   4
CH3COHCH3               C   3H   7O   1     G    300.00   4000.00 1388.00      1
 .115026438E+02 .149881248E-01-.510421075E-05 .789864272E-09-.457135659E-13    2
-.164821894E+05-.347655748E+02 .118802517E+01 .410410262E-01-.314650841E-04    3
 .133514692E-07-.237788249E-11-.130177234E+05 .200655998E+02                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   4000.00 1674.00      1
 .931287816E+01 .167579212E-01-.575555480E-05 .900584362E-09-.526566836E-13    2
-.119163093E+05-.195564662E+02 .120494302E+01 .330857885E-01-.163893637E-04    3
 .318103918E-08-.684229288E-13-.902896295E+04 .246601603E+02                   4
CH3CO2H                 C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .767084601E+01 .135152602E-01-.525874333E-05 .893184479E-09-.553180543E-13    2
-.557560970E+05-.154677315E+02 .278950201E+01 .999941719E-02 .342572245E-04    3
-.509031329E-07 .206222185E-10-.534752488E+05 .141053123E+02                   4
HCOOH                   C   1H   2O   2     G    300.00   4000.00 1000.00      1        POLIMI
 .461383160E+01 .644963640E-02-.229082510E-05 .367160470E-09-.218736750E-13    2
-.453303180E+05 .847883830E+00 .389836160E+01-.355877950E-02 .355205380E-04    3
-.438499590E-07 .171077690E-10-.467785744E+05 .734953970E+01                   4
HCO3                    C   1H   1O   3     G    300.00   4000.00 1000.00      1
 .726425669E+01 .532196974E-02-.196520055E-05 .323182996E-09-.195989250E-13    2
-.159242239E+05-.103647520E+02 .364808935E+01 .957717212E-02 .755287366E-05    3
-.181264650E-07 .827293980E-11-.146544449E+05 .967735548E+01                   4
HCO3H                   C   1H   2O   3     G    300.00   4000.00 1378.00      1
 .987503581E+01 .464663708E-02-.167230522E-05 .268624413E-09-.159595232E-13    2
-.380502456E+05-.224938942E+02 .242464726E+01 .219706380E-01-.168705546E-04    3
 .625612194E-08-.911645843E-12-.354828006E+05 .175027796E+02                   4
H2                TPIS78H   2    0    0    0G   200.000  6000.00  1000.00      1
 2.93286575E+00 8.26608026E-04-1.46402364E-07 1.54100414E-11-6.88804800E-16    2
-8.13065581E+02-1.02432865E+00 2.34433112E+00 7.98052075E-03-1.94781510E-05    3
 2.01572094E-08-7.37611761E-12-9.17935173E+02 6.83010238E-01 0.00000000E+00    4
H                 L 6/94H   1    0    0    0G   200.000  6000.00  1000.00      1
 0.25000000E+01 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.25473660E+05-0.44668285E+00 0.25000000E+01 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.25473660E+05-0.44668285E+00 0.26219035E+05    4
O2                RUS 89O   2    0    0    0G   200.000  6000.00  1000.00      1
 3.66096065E+00 6.56365811E-04-1.41149627E-07 2.05797935E-11-1.29913436E-15    2
-1.21597718E+03 3.41536279E+00 3.78245636E+00-2.99673416E-03 9.84730201E-06    3
-9.68129509E-09 3.24372837E-12-1.06394356E+03 3.65767573E+00 0.00000000E+00    4
O                 L 1/90O   1    0    0    0G   200.000  6000.00  1000.00      1
 2.54363697E+00-2.73162486E-05-4.19029520E-09 4.95481845E-12-4.79553694E-16    2
 2.92260120E+04 4.92229457E+00 3.16826710E+00-3.27931884E-03 6.64306396E-06    3
-6.12806624E-09 2.11265971E-12 2.91222592E+04 2.05193346E+00 2.99687009E+04    4
H2O               L 5/89H   2 O  1    0    0G   200.000  6000.00  1000.00      1
 0.26770389E+01 0.29731816E-02-0.77376889E-06 0.94433514E-10-0.42689991E-14    2
-0.29885894E+05 0.68825500E+01 0.41986352E+01-0.20364017E-02 0.65203416E-05    3
-0.54879269E-08 0.17719680E-11-0.30293726E+05-0.84900901E+00-0.29084817E+05    4
OH                IU3/03O   1 H  1    0    0G   200.000  6000.00  1000.00      1
 2.83853033E+00 1.10741289E-03-2.94000209E-07 4.20698729E-11-2.42289890E-15    2
 3.69780808E+03 5.84494652E+00 3.99198424E+00-2.40106655E-03 4.61664033E-06    3
-3.87916306E-09 1.36319502E-12 3.36889836E+03-1.03998477E-01 4.48613328E+03    4
OHV               121286O   1H   1          G  0300.00   5000.00  1000.00      1
 0.02882730E+02 0.10139743E-02-0.02276877E-05 0.02174683E-09-0.05126305E-14    2
 5.02650000E+04 0.05595712E+02 0.03637266E+02 0.01850910E-02-0.16761646E-05    3
 0.02387202E-07-0.08431442E-11 5.00213000E+04 0.13588605E+01                   4
H2O2              T 8/03H   2O   2    0    0G   200.000  6000.00  1000.00      1
 4.57977305E+00 4.05326003E-03-1.29844730E-06 1.98211400E-10-1.13968792E-14    2
-1.80071775E+04 6.64970694E-01 4.31515149E+00-8.47390622E-04 1.76404323E-05    3
-2.26762944E-08 9.08950158E-12-1.77067437E+04 3.27373319E+00-1.63425145E+04    4
HO2               T 1/09H   1O   2    0    0G   200.000  5000.00  1000.00      1
 4.17228741E+00 1.88117627E-03-3.46277286E-07 1.94657549E-11 1.76256905E-16    2
 3.10206839E+01 2.95767672E+00 4.30179807E+00-4.74912097E-03 2.11582905E-05    3
-2.42763914E-08 9.29225225E-12 2.64018485E+02 3.71666220E+00 1.47886045E+03    4
CO                RUS 79C   1O   1    0    0G   200.000  6000.00  1000.00      1
 0.30484859E+01 0.13517281E-02-0.48579405E-06 0.78853644E-10-0.46980746E-14    2
-0.14266117E+05 0.60170977E+01 0.35795335E+01-0.61035369E-03 0.10168143E-05    3
 0.90700586E-09-0.90442449E-12-0.14344086E+05 0.35084093E+01-0.13293628E+05    4
CO2               L 7/88C   1O   2    0    0G   200.000  6000.00  1000.00      1
 0.46365111E+01 0.27414569E-02-0.99589759E-06 0.16038666E-09-0.91619857E-14    2
-0.49024904E+05-0.19348955E+01 0.23568130E+01 0.89841299E-02-0.71220632E-05    3
 0.24573008E-08-0.14288548E-12-0.48371971E+05 0.99009035E+01-0.47328105E+05    4
HOCO              T05/06H  1 C  1 O  2    0 G   200.000  6000.00   1000.00     1
 5.39206152E+00 4.11221455E-03-1.48194900E-06 2.39875460E-10-1.43903104E-14    2
-2.38606717E+04-2.23529091E+00 2.92207919E+00 7.62453859E-03 3.29884437E-06    3
-1.07135205E-08 5.11587057E-12-2.30281524E+04 1.12925886E+01-2.18076591E+04    4
CH4               G 8/99C  1 H  4    0    0 G   200.000  6000.00  1000.00      1
 1.65326226E+00 1.00263099E-02-3.31661238E-06 5.36483138E-10-3.14696758E-14    2
-1.00095936E+04 9.90506283E+00 5.14911468E+00-1.36622009E-02 4.91453921E-05    3
-4.84246767E-08 1.66603441E-11-1.02465983E+04-4.63848842E+00-8.97226656E+03    4
CH3               IU0702C  1 H  3    0    0 G   200.000  6000.00  1000.00      1
 0.29781206E+01 0.57978520E-02-0.19755800E-05 0.30729790E-09-0.17917416E-13    2
 0.16509513E+05 0.47224799E+01 0.36571797E+01 0.21265979E-02 0.54583883E-05    3
-0.66181003E-08 0.24657074E-11 0.16422716E+05 0.16735354E+01 0.17643935E+05    4
CH2               IU3/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
 3.14631886E+00 3.03671259E-03-9.96474439E-07 1.50483580E-10-8.57335515E-15    2
 4.60412605E+04 4.72341711E+00 3.71757846E+00 1.27391260E-03 2.17347251E-06    3
-3.48858500E-09 1.65208866E-12 4.58723866E+04 1.75297945E+00 4.70504920E+04    4
CH2(S)            IU6/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
 3.13501686E+00 2.89593926E-03-8.16668090E-07 1.13572697E-10-6.36262835E-15    2
 5.05040504E+04 4.06030621E+00 4.19331325E+00-2.33105184E-03 8.15676451E-06    3
-6.62985981E-09 1.93233199E-12 5.03662246E+04-7.46734310E-01 5.15727280E+04    4
C                 L 7/88C   1     0    0   0G   200.000  6000.00  1000.00      1
 0.26055830E+01-0.19593434E-03 0.10673722E-06-0.16423940E-10 0.81870580E-15    2
 0.85411742E+05 0.41923868E+01 0.25542395E+01-0.32153772E-03 0.73379223E-06    3
-0.73223487E-09 0.26652144E-12 0.85442681E+05 0.45313085E+01 0.86195097E+05    4
CH                IU3/03C  1 H  1    0    0 G   200.000  6000.00  1000.00      1
 0.25209369E+01 0.17653639E-02-0.46147660E-06 0.59289675E-10-0.33474501E-14    2
 0.70946769E+05 0.74051829E+01 0.34897583E+01 0.32432160E-03-0.16899751E-05    3
 0.31628420E-08-0.14061803E-11 0.70612646E+05 0.20842841E+01 0.71658188E+05    4
CHV               073003C   1H   1          G  0300.00   5000.00  1000.00      1
 0.02196223E+02 0.02340381E-01-0.07058201E-05 0.09007582E-09-0.03855040E-13    2
 0.10419559E+06 0.09178373E+02 0.03200202E+02 0.02072875E-01-0.05134431E-04    3
 0.05733890E-07-0.01955533E-10 0.10393714E+06 0.03331587E+02                   4
CH3O2H            A 7/05C  1 H  4 O  2    0 G   200.000  6000.00  1000.00      1
 7.76538058E+00 8.61499712E-03-2.98006935E-06 4.68638071E-10-2.75339255E-14    2
-1.82979984E+04-1.43992663E+01 2.90540897E+00 1.74994735E-02 5.28243630E-06    3
-2.52827275E-08 1.34368212E-11-1.68894632E+04 1.13741987E+01-1.52423685E+04    4
CH3O2                   H   3C   1O   2    0G   300.000  5000.000 1374.000    11
 6.47970487E+00 7.44401080E-03-2.52348555E-06 3.89577296E-10-2.25182399E-14    2
-1.56285441E+03-8.19477074E+00 1.97339205E+00 1.53542340E-02-6.37314891E-06    3
 3.19930565E-10 2.82193915E-13 2.54278835E+02 1.69194215E+01                   4
CH2O2H     9/ 1/12      C   1H   3O   2    0G   300.000  5000.000 1410.000    21
 9.24697852E+00 4.60845541E-03-1.53501472E-06 2.34434830E-10-1.34573106E-14    2
 4.11529953E+03-2.11503248E+01 2.88976454E+00 2.09465776E-02-1.75190772E-05    3
 7.27819787E-09-1.18912344E-12 6.12390620E+03 1.23802076E+01                   4
CH3OH             T06/02C   1H  4 O  1    0 G   200.000  6000.00  1000.00      1
 3.52726795E+00 1.03178783E-02-3.62892944E-06 5.77448016E-10-3.42182632E-14    2
-2.60028834E+04 5.16758693E+00 5.65851051E+00-1.62983419E-02 6.91938156E-05    3
-7.58372926E-08 2.80427550E-11-2.56119736E+04-8.97330508E-01-2.41746056E+04    4
CH3O              IU1/03C  1 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 4.75779238E+00 7.44142474E-03-2.69705176E-06 4.38090504E-10-2.63537098E-14    2
 3.78111940E+02-1.96680028E+00 3.71180502E+00-2.80463306E-03 3.76550971E-05    3
-4.73072089E-08 1.86588420E-11 1.29569760E+03 6.57240864E+00 2.52571660E+03    4
CH2OH             IU2/03C  1 H  3 O  1    0 G   200.000  6000.00   1000.00     1
 5.09314370E+00 5.94761260E-03-2.06497460E-06 3.23008173E-10-1.88125902E-14    2
-4.03409640E+03-1.84691493E+00 4.47834367E+00-1.35070310E-03 2.78484980E-05    3
-3.64869060E-08 1.47907450E-11-3.50072890E+03 3.30913500E+00-2.04462770E+03    4
CH2O              T 5/11H   2C   1O   1    0G   200.000  6000.00  1000.00      1
 3.16952665E+00 6.19320560E-03-2.25056366E-06 3.65975660E-10-2.20149458E-14    2
-1.45486831E+04 6.04207898E+00 4.79372312E+00-9.90833322E-03 3.73219990E-05    3
-3.79285237E-08 1.31772641E-11-1.43791953E+04 6.02798058E-01-1.31293365E+04    4
HCO               T 5/03C  1 H  1 O  1    0 G   200.000  6000.00  1000.00      1
 3.92001542E+00 2.52279324E-03-6.71004164E-07 1.05615948E-10-7.43798261E-15    2
 3.65342928E+03 3.58077056E+00 4.23754610E+00-3.32075257E-03 1.40030264E-05    3
-1.34239995E-08 4.37416208E-12 3.87241185E+03 3.30834869E+00 5.08749163E+03    4
HCOH              MAR94 C   1H   2O   1    0G   300.     5000.    1398.        1
 9.18749272E+00 1.52011152E-03-6.27603516E-07 1.09727989E-10-6.89655128E-15    2
 7.81364593E+03-2.73434214E+01-2.82157421E+00 3.57331702E-02-3.80861580E-05    3
 1.86205951E-08-3.45957838E-12 1.12956672E+04 3.48487757E+01                   4
HO2CHO     6/26/95 THERMC   1H   2O   3    0G   300.000  5000.000 1378.00     21
 9.87503878E+00 4.64663708E-03-1.67230522E-06 2.68624413E-10-1.59595232E-14    2
-3.80502496E+04-2.24939155E+01 2.42464726E+00 2.19706380E-02-1.68705546E-05    3
 6.25612194E-09-9.11645843E-13-3.54828006E+04 1.75027796E+01                   4
HOCH2O2H   9/ 1/12      C   1H   4O   3    0G   300.000  5000.000 1398.000    21
 1.24531886E+01 7.18221110E-03-2.47029548E-06 3.85611737E-10-2.24774193E-14    2
-4.24862928E+04-3.58745197E+01 5.35189713E-01 3.73266553E-02-3.15299511E-05    3
 1.30352583E-08-2.11473264E-12-3.86609415E+04 2.71776082E+01                   4
HOCH2O2    9/ 1/12      C   1H   3O   3    0G   300.000  5000.000 1377.000    21
 1.16406115E+01 5.72826040E-03-2.05362036E-06 3.29070695E-10-1.95188360E-14    2
-2.53505769E+04-3.07332064E+01 2.82068616E+00 2.47857094E-02-1.66186399E-05    3
 4.79633095E-09-4.28087766E-13-2.22077036E+04 1.70599803E+01                   4
OCH2O2H    7/21/14 THERMC   1H   3O   3    0G   300.000  5000.000 1418.000    31
 1.29622491E+01 4.21948855E-03-1.54275194E-06 2.50413077E-10-1.49855537E-14    2
-1.81326406E+04-3.87016356E+01 4.46349361E-01 3.63049606E-02-3.26130978E-05    3
 1.37050551E-08-2.20872791E-12-1.41972598E+04 2.72960376E+01                   4
HOCH2O     2/16/99 THERMC   1H   3O   2    0G   300.000  5000.000 1452.000    11
 6.39521515E+00 7.43673043E-03-2.50422354E-06 3.84879712E-10-2.21778689E-14    2
-2.41108840E+04-6.63865583E+00 4.11183145E+00 7.53850697E-03 3.77337370E-06    3
-5.38746005E-09 1.45615887E-12-2.28023001E+04 7.46807254E+00                   4
O2CHO      6/26/95 THERMC   1H   1O   3    0G   300.000  5000.000 1368.00     11
 7.24075139E+00 4.63312951E-03-1.63693995E-06 2.59706693E-10-1.52964699E-14    2
-1.87027618E+04-6.49547212E+00 3.96059309E+00 1.06002279E-02-5.25713351E-06    3
 1.01716726E-09-2.87487602E-14-1.73599383E+04 1.17807483E+01                   4
HOCHO             L 8/88H   2C   1O   2    0G   200.000  6000.00  1000.00      1
 0.46138316E+01 0.64496364E-02-0.22908251E-05 0.36716047E-09-0.21873675E-13    2
-0.47514850E+05 0.84788383E+00 0.38983616E+01-0.35587795E-02 0.35520538E-04    3
-0.43849959E-07 0.17107769E-10-0.46770609E+05 0.73495397E+01-0.45531246E+05    4
OCHO              ATCT/AC  1 O  2 H  1    0 G   200.000  6000.000 1000.00      1
 4.14394211E+00 5.59738818E-03-1.99794019E-06 3.16179193E-10-1.85614483E-14    2
-1.72459887E+04 5.07778617E+00 4.68825921E+00-4.14871834E-03 2.55066010E-05    3
-2.84473900E-08 1.04422559E-11-1.69867041E+04 4.28426480E+00-1.55992356E+04    4
C2H6              G 8/88C   2H 6    0      0G   200.000  6000.00  1000.00      1
 4.04666411E+00 1.53538802E-02-5.47039485E-06 8.77826544E-10-5.23167531E-14    2
-1.24473499E+04-9.68698313E-01 4.29142572E+00-5.50154901E-03 5.99438458E-05    3
-7.08466469E-08 2.68685836E-11-1.15222056E+04 2.66678994E+00-1.00849652E+04    4
C2H5       8/ 4/ 4 THERMC   2H   5    0    0G   300.000  5000.000 1387.000    11
 5.88784390E+00 1.03076793E-02-3.46844396E-06 5.32499257E-10-3.06512651E-14    2
 1.15065499E+04-8.49651771E+00 1.32730217E+00 1.76656753E-02-6.14926558E-06    3
-3.01143466E-10 4.38617775E-13 1.34284028E+04 1.71789216E+01                   4
C2H5O2H    9/ 1/12      C   2H   6O   2    0G   300.000  5000.000 1390.000    31
 1.04823538E+01 1.34779879E-02-4.62179078E-06 7.18618519E-10-4.17307436E-14    2
-2.46578171E+04-2.84294243E+01 1.83755328E+00 3.38053586E-02-2.37548140E-05    3
 9.31974865E-09-1.58003428E-12-2.15814086E+04 1.80977584E+01                   4
C2H5O2     9/ 1/12      C   2H   5O   2    0G   300.000  5000.000 1389.000    21
 9.50282570E+00 1.20429839E-02-4.09491581E-06 6.33049241E-10-3.66133788E-14    2
-7.37069391E+03-2.21717130E+01 3.90351912E+00 2.22599212E-02-1.01610079E-05    3
 1.71709751E-09 1.88166738E-14-5.09654081E+03 8.98722750E+00                   4
C2H4       8/12/15      C   2H   4    0    0G   300.000  5000.000 1392.000    01
 5.07061289E+00 9.11140768E-03-3.10506692E-06 4.80733851E-10-2.78321396E-14    2
 3.66391217E+03-6.64501414E+00 4.81118223E-01 1.83778060E-02-9.99633565E-06    3
 2.73211039E-09-3.01837289E-13 5.44386648E+03 1.85867157E+01                   4
C2H3       8/12/15      C   2H   3    0    0G   300.000  5000.000 1400.000    01
 4.99675415E+00 6.55838271E-03-2.20921909E-06 3.39300272E-10-1.95316926E-14    2
 3.34604382E+04-3.01451097E+00 1.25545094E+00 1.57481597E-02-1.12218328E-05    3
 4.50915682E-09-7.74861577E-13 3.47435574E+04 1.69664043E+01                   4
CHOCHO                  C   2H   2O   2    0G   300.000  5000.000 1386.000    11
 9.75438561E+00 4.97645947E-03-1.74410483E-06 2.75586994E-10-1.61969892E-14    2
-2.95832896E+04-2.61878329E+01 1.88105120E+00 2.36386368E-02-1.83443295E-05    3
 6.84842963E-09-9.92733674E-13-2.69280190E+04 1.59154793E+01                   4
C2H3OOH    4/18/ 8 THERMC   2H   4O   2    0G   300.000  5000.000 1397.000    21
 1.15749951E+01 8.09909174E-03-2.81808668E-06 4.42697954E-10-2.58998042E-14    2
-8.84852664E+03-3.43859117E+01 1.35644398E+00 3.37002447E-02-2.75988500E-05    3
 1.14222854E-08-1.89488886E-12-5.49996692E+03 1.98354466E+01                   4
C2H3OO                  H   3C   2O   2     G   298.150  2000.000 1000.00      1
 6.04483828E+00 1.45511127E-02-7.50974622E-06 1.83488280E-09-1.66689681E-13    2
 1.01699244E+04-3.71144913E+00 1.09784776E+00 2.95333237E-02-2.27744360E-05    3
 7.20559155E-09-3.07929092E-13 1.13996101E+04 2.13563583E+01                   4
CHCHO                   H   2C   2O   1     G   298.150  2000.000 1000.00      1
 4.92632910E+00 9.71712147E-03-5.54855980E-06 1.53068537E-09-1.64742462E-13    2
 2.89499494E+04 5.27874677E-01 2.33256751E+00 1.62952986E-02-9.72052177E-06    3
 5.15124155E-10 1.03836514E-12 2.96585452E+04 1.39904923E+01                   4
C2H2              G 1/91C  2 H  2    0    0 G   200.000  6000.00  1000.00      1
 4.65878489E+00 4.88396667E-03-1.60828888E-06 2.46974544E-10-1.38605959E-14    2
 2.57594042E+04-3.99838194E+00 8.08679682E-01 2.33615762E-02-3.55172234E-05    3
 2.80152958E-08-8.50075165E-12 2.64289808E+04 1.39396761E+01 2.74459950E+04    4
C2H               T 5/10C  2 H  1    0    0 G   200.000  6000.00  1000.00      1
 3.66270248E+00 3.82492252E-03-1.36632500E-06 2.13455040E-10-1.23216848E-14    2
 6.71683790E+04 3.92205792E+00 2.89867676E+00 1.32988489E-02-2.80733327E-05    3
 2.89484755E-08-1.07502351E-11 6.70616050E+04 6.18547632E+00 6.83210436E+04    4
H2CC              L12/89H   2C   2    0    0G   200.000  6000.000  1000.000    1
 0.42780340E+01 0.47562804E-02-0.16301009E-05 0.25462806E-09-0.14886379E-13    2
 0.48316688E+05 0.64023701E+00 0.32815483E+01 0.69764791E-02-0.23855244E-05    3
-0.12104432E-08 0.98189545E-12 0.48621794E+05 0.59203910E+01 0.49887266E+05    4
C2H5OH     8/12/15      C   2H   6O   1    0G   300.000  5000.000 1402.000    21
 8.14483865E+00 1.28314052E-02-4.29052743E-06 6.55971721E-10-3.76506611E-14    2
-3.24005526E+04-1.86241126E+01 2.15805861E-01 2.95228396E-02-1.68271048E-05    3
 4.49484797E-09-4.02451543E-13-2.94851823E+04 2.45725052E+01                   4
C2H5O      8/12/15      C   2H   5O   1    0G   300.000  5000.000 1467.000    11
 8.19120635E+00 1.10391986E-02-3.75270536E-06 5.80275784E-10-3.35735146E-14    2
-5.66847208E+03-1.90131344E+01 2.90353584E+00 1.77256708E-02-2.69624757E-06    3
-3.45830533E-09 1.25224784E-12-3.28930290E+03 1.13545591E+01                   4
PC2H4OH    8/12/15      C   2H   5O   1    0G   300.000  5000.000 1395.000    21
 8.06750150E+00 1.06143554E-02-3.57999360E-06 5.50363760E-10-3.17051769E-14    2
-6.92747939E+03-1.53833428E+01 2.59479867E+00 2.27100669E-02-1.39473846E-05    3
 4.70095591E-09-6.90044236E-13-4.91486975E+03 1.43240718E+01                   4
SC2H4OH    8/12/15      C   2H   5O   1    0G   300.000  5000.000 1385.000    21
 8.15007136E+00 1.02549305E-02-3.40137764E-06 5.17509965E-10-2.96128942E-14    2
-1.05014386E+04-1.73134615E+01 1.46281093E+00 2.39193995E-02-1.30667185E-05    3
 3.10615465E-09-1.85896007E-13-8.00790323E+03 1.92547092E+01                   4
O2C2H4OH   9/ 1/12 THERMC   2H   5O   3    0G   300.000  5000.000 1506.000    41
 1.27503881E+01 1.11514325E-02-3.83473891E-06 5.98155829E-10-3.48372108E-14    2
-2.52770876E+04-3.54317608E+01 7.04009800E+00 1.59564166E-02 2.21097416E-06    3
-7.05197355E-09 2.08266026E-12-2.24524432E+04-1.75361758E+00                   4
C2H4O2H    9/ 1/12      C   2H   5O   2    0G   300.000  5000.000 1389.000    31
 1.00590614E+01 1.13378955E-02-3.89403387E-06 6.06090687E-10-3.52212353E-14    2
 4.24048653E+02-2.32086536E+01 2.75788364E+00 2.88271987E-02-2.08302264E-05    3
 8.47401397E-09-1.48617610E-12 3.00153893E+03 1.59921711E+01                   4
C2H4O1-2          L 8/88C  2 H  4 O  1    0 G   200.000  6000.00  1000.00      1
 0.54887641E+01 0.12046190E-01-0.43336931E-05 0.70028311E-09-0.41949088E-13    2
-0.91804251E+04-0.70799605E+01 0.37590532E+01-0.94412180E-02 0.80309721E-04    3
-0.10080788E-06 0.40039921E-10-0.75608143E+04 0.78497475E+01-0.63304657E+04    4
C2H3O1-2          A 1/05C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 5.60158035E+00 9.17613962E-03-3.28028902E-06 5.27903888E-10-3.15362241E-14    2
 1.71446252E+04-5.47228512E+00 3.58349017E+00-6.02275805E-03 6.32426867E-05    3
-8.18540707E-08 3.30444505E-11 1.85681353E+04 9.59725926E+00 1.97814471E+04    4
CH3CHO            L 8/88C  2 H  4 O   1   0 G   200.000  6000.00  1000.00      1
 0.54041108E+01 0.11723059E-01-0.42263137E-05 0.68372451E-09-0.40984863E-13    2
-0.22593122E+05-0.34807917E+01 0.47294595E+01-0.31932858E-02 0.47534921E-04    3
-0.57458611E-07 0.21931112E-10-0.21572878E+05 0.41030159E+01-0.19987949E+05    4
CH3CO             IU2/03C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 0.53137165E+01 0.91737793E-02-0.33220386E-05 0.53947456E-09-0.32452368E-13    2
-0.36450414E+04-0.16757558E+01 0.40358705E+01 0.87729487E-03 0.30710010E-04    3
-0.39247565E-07 0.15296869E-10-0.26820738E+04 0.78617682E+01-0.12388039E+04    4
CH2CHO            T03/10C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 6.53928338E+00 7.80238629E-03-2.76413612E-06 4.42098906E-10-2.62954290E-14    2
-1.18858659E+03-8.72091393E+00 2.79502600E+00 1.01099472E-02 1.61750645E-05    3
-3.10303145E-08 1.39436139E-11 1.62944975E+02 1.23646657E+01 1.53380440E+03    4
O2CH2CHO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1393.000    01
 1.11807543E+01 9.14479256E-03-3.15089833E-06 4.91944238E-10-2.86639180E-14    2
-1.55790331E+04-2.87892740E+01-1.29465843E+00 4.44936393E-02-4.26577074E-05    3
 2.07391950E-08-3.96828771E-12-1.18275628E+04 3.60778797E+01                   4
HO2CH2CO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1386.000    01
 1.04146322E+01 1.12680116E-02-5.17494839E-06 1.00333285E-09-6.68165911E-14    2
-1.40955672E+04-2.27894400E+01 2.22681686E+00 3.56781380E-02-3.26401909E-05    3
 1.47651988E-08-2.64794380E-12-1.18735095E+04 1.91581197E+01                   4
C2H3OH     2/ 3/ 9 THERMC   2H   4O   1    0G   300.000  5000.000 1410.000    11
 8.32598158E+00 8.03387281E-03-2.63928405E-06 3.98410726E-10-2.26551155E-14    2
-1.83221436E+04-2.02080305E+01-1.27972260E-01 3.38506073E-02-3.30644935E-05    3
 1.64858739E-08-3.19935455E-12-1.59914544E+04 2.30438601E+01                   4
C2H2OH                  H   3C   2O   1    0G   300.000  5000.000 1401.000    11
 8.20268447E+00 5.92989165E-03-1.99194448E-06 3.05794341E-10-1.76114732E-14    2
 1.24881328E+04-1.89670436E+01 6.41642616E-01 2.61903633E-02-2.30385370E-05    3
 1.02804704E-08-1.81971416E-12 1.48276951E+04 2.06750999E+01                   4
CH2CO                   H   2C   2O   1    0G    300.00   5000.00 1000.00      1
 5.35869367E+00 6.95641586E-03-2.64802637E-06 4.65067592E-10-3.08641820E-14    2
-7.90294013E+03-3.98525731E+00 1.81422511E+00 1.99008590E-02-2.21416008E-05    3
 1.45028521E-08-3.98877068E-12-7.05394926E+03 1.36079359E+01                   4
HCCO              T 4/09H  1 C  2 O  1    0 G   200.000  6000.00  1000.00      1
 5.91479333E+00 3.71408730E-03-1.30137010E-06 2.06473345E-10-1.21476759E-14    2
 1.93596301E+04-5.50567269E+00 1.87607969E+00 2.21205418E-02-3.58869325E-05    3
 3.05402541E-08-1.01281069E-11 2.01633840E+04 1.36968290E+01 2.14444387E+04    4
HCCOH             T12/09C  2 H  2 O  1    0 G   200.000  6000.00  1000.00      1
 6.37509678E+00 5.49429011E-03-1.88136576E-06 2.93803536E-10-1.71771901E-14    2
 8.93277676E+03-8.24498007E+00 2.05541154E+00 2.52003372E-02-3.80821654E-05    3
 3.09890632E-08-9.89799902E-12 9.76872113E+03 1.22271534E+01 1.12217316E+04    4
CH3CO3H    6/26/95 THERMC   2H   4O   3    0G   300.000  5000.000 1391.000    31
 1.25060485E+01 9.47789695E-03-3.30402246E-06 5.19630793E-10-3.04233568E-14    2
-4.59856703E+04-3.79195947E+01 2.24135876E+00 3.37963514E-02-2.53887482E-05    3
 9.67583587E-09-1.49266157E-12-4.24677831E+04 1.70668133E+01                   4
CH3CO3     4/ 3/ 0 THERMC   2H   3O   3    0G   300.000  5000.000 1391.000    21
 1.12522498E+01 8.33652672E-03-2.89014530E-06 4.52781734E-10-2.64354456E-14    2
-2.60238584E+04-2.96370457E+01 3.60373432E+00 2.70080341E-02-2.08293438E-05    3
 8.50541104E-09-1.43846110E-12-2.34205171E+04 1.12014914E+01                   4
CH3CO2     2/14/95 THERMC   2H   3O   2    0G   300.000  5000.000 1395.000    11
 8.54059736E+00 8.32951214E-03-2.84722010E-06 4.41927196E-10-2.56373394E-14    2
-2.97290678E+04-2.03883545E+01 1.37440768E+00 2.49115604E-02-1.74308894E-05    3
 6.24799508E-09-9.09516835E-13-2.72330150E+04 1.81405454E+01                   4
!CH3OCH3    2/11/14 THERMC   2H   6O   1    0G   300.000  5000.000 1999.000    21
! 6.03232751E+00 1.56155270E-02-5.50761030E-06 8.75666140E-10-5.17180562E-14    2
!-2.52690354E+04-8.25885183E+00 2.05597390E+00 2.07019456E-02-5.00382376E-06    3
!-1.62279885E-09 6.84330155E-13-2.35494445E+04 1.45029944E+01                   4
!CH3OCH2    2/11/14 THERMC   2H   5O   1    0G   300.000  5000.000 1395.000    11
! 6.62621974E+00 1.22219496E-02-4.12416696E-06 6.34127512E-10-3.65317390E-14    2
!-3.33965890E+03-8.95305753E+00 1.58874948E+00 2.24414123E-02-1.19434933E-05    3
! 3.37160213E-09-4.15077249E-13-1.37208255E+03 1.87548958E+01                   4
CHOCHO                  C   2H   2O   2     G    300.00   4000.00 1000.00      1
 .872506895E+01 .633096819E-02-.235574814E-05 .389782853E-09-.237486912E-13    2
-.291024131E+05-.203903909E+02 .468412461E+01 .478012819E-03 .426390768E-04    3
-.579018239E-07 .231669328E-10-.271985007E+05 .451187184E+01                   4
CH2OHCHO                C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .691088832E+01 .123280849E-01-.438373062E-05 .703055164E-09-.419009846E-13    2
-.400211587E+05-.696132551E+01 .614926095E+01-.596828114E-02 .596003337E-04    3
-.716663578E-07 .274014411E-10-.388356849E+05 .186644598E+01                   4
O2C2H4O2H               C   2H   5O   4     G    300.00   4000.00 1387.00      1
 .145471032E+02 .123393823E-01-.427259469E-05 .668763337E-09-.390196721E-13    2
-.196338761E+05-.408784236E+02 .590031872E+01 .305658528E-01-.185905950E-04    3
 .567871605E-08-.702799577E-12-.163916571E+05 .633051038E+01                   4
HO2CH2CHO               C   2H   4O   3     G    300.00   4000.00 1000.00      1
 .127662941E+02 .102143437E-01-.363547001E-05 .583491588E-09-.347179974E-13    2
-.753528536E+05-.396511752E+02 .280443702E+01 .210851644E-01 .335863233E-04    3
-.702669107E-07 .326849274E-10-.720649998E+05 .151180675E+02                   4
CH3OCH2O2H 2/12/14 THERMC   2H   6O   3    0G   300.000  5000.000 1404.000    31
 1.28159161E+01 1.34818095E-02-4.50397729E-06 6.88229286E-10-3.94883680E-14    2
-4.06745921E+04-3.78047802E+01 1.05786981E+00 4.36787095E-02-3.46383899E-05    3
 1.44808830E-08-2.46100643E-12-3.68851076E+04 2.43391936E+01                   4
CH3OCH2O2  2/12/14 THERMC   2H   5O   3    0G   300.000  5000.000 1441.000    21
 1.19179361E+01 1.19412867E-02-3.93526185E-06 5.95756132E-10-3.39597705E-14    2
-2.34231833E+04-3.20096863E+01 3.39930541E+00 3.09460407E-02-1.92548181E-05    3
 5.76033887E-09-6.16081571E-13-2.04433218E+04 1.39429608E+01                   4
CH2OCH2O2H 2/12/14 THERMC   2H   5O   3    0G   300.000  5000.000 1418.000    21
 1.23892901E+01 1.11758961E-02-3.59249095E-06 5.34196366E-10-3.00536541E-14    2
-1.80551598E+04-3.29576862E+01 1.62245477E-01 4.76101093E-02-4.52046954E-05    3
 2.18379311E-08-4.11295947E-12-1.46498100E+04 2.98253164E+01                   4
O2CH2OCH2O2H 2/12/14 ERMC   2H   5O   5    0G   300.000  5000.000 1433.000    31
 1.77378326E+01 1.13589899E-02-3.67382539E-06 5.49255712E-10-3.10405899E-14    2
-3.82903058E+04-5.66609932E+01 2.39977678E+00 5.39881943E-02-4.87969524E-05    3
 2.19792134E-08-3.86106979E-12-3.37824638E+04 2.30683371E+01                   4
HO2CH2OCHO 2/12/14 THERMC   2H   4O   4    0G   300.000  5000.000 1386.000    31
 1.57136128E+01 9.64430166E-03-3.44136025E-06 5.49722196E-10-3.25360322E-14    2
-6.29409094E+04-5.29505242E+01 1.21909586E+00 4.28858235E-02-3.17634222E-05    3
 1.11542676E-08-1.49753153E-12-5.79287926E+04 2.49759193E+01                   4
OCH2OCHO   5/29/14 THERMC   2H   3O   3    0G   300.000  5000.000 1523.000    21
 1.24013200E+01 7.83738243E-03-2.82992688E-06 4.55558739E-10-2.71061389E-14    2
-4.68453470E+04-3.78084549E+01 1.89539692E+00 2.74118545E-02-1.36476090E-05    3
 1.26325603E-09 5.17970476E-13-4.27879440E+04 2.02333278E+01                   4
HOCH2OCO   5/29/14 THERMC   2H   3O   3    0G   300.000  5000.000 1443.000    11
 1.11498410E+01 9.34736520E-03-3.35541548E-06 5.38037115E-10-3.19260183E-14    2
-4.75012119E+04-2.95983867E+01 5.95255071E+00 8.42196282E-03 1.36741678E-05    3
-1.46786275E-08 3.84143533E-12-4.44470269E+04 2.85657217E+00                   4
CH3OCH2O   5/15/14 THERMC   2H   5O   2    0G   300.000  5000.000 1523.000    31
 9.81288609E+00 1.21313106E-02-4.30285768E-06 6.84443177E-10-4.03862658E-14    2
-2.50760742E+04-2.51866352E+01 5.63414373E+00 8.92830283E-03 1.37225633E-05    3
-1.40497059E-08 3.54625624E-12-2.22825214E+04 1.93588846E+00                   4
CH3OCHO           T 6/08C  2 H  4 O  2    0 G   200.000  6000.00  1000.00      1
 6.33360880E+00 1.34851485E-02-4.84305805E-06 7.81719241E-10-4.67917447E-14    2
-4.68316521E+04-6.91542601E+00 5.96757028E+00-9.38085425E-03 7.07648417E-05    3
-8.29932227E-08 3.13522917E-11-4.55713267E+04 7.50341113E-01-4.37330508E+04    4
CH3OCO     5/ 8/ 3 THERMC   2H   3O   2    0G   300.000  5000.000 1601.000    21
 9.73659803E+00 7.42432713E-03-2.65641779E-06 4.25031143E-10-2.51824924E-14    2
-2.36015721E+04-2.36353471E+01 4.16215406E+00 1.38037511E-02-3.08486109E-07    3
-4.56430814E-09 1.46909632E-12-2.10130301E+04 8.64301044E+00                   4
CH2OCHO    4/15/ 8 THERMC   2H   3O   2    0G   300.000  5000.000 1442.000    21
 1.00960096E+01 7.19887066E-03-2.59813465E-06 4.18110812E-10-2.48723387E-14    2
-2.36389018E+04-2.71144175E+01 2.31031671E+00 1.80474065E-02-2.71519637E-06    3
-4.60918579E-09 1.70037078E-12-2.02910878E+04 1.71549722E+01                   4
C3H8       8/12/15      C   3H   8    0    0G   300.000  5000.000 1390.000    21
 9.15541310E+00 1.72574139E-02-5.85614868E-06 9.04190155E-10-5.22523772E-14    2
-1.75762439E+04-2.77418510E+01 2.40878470E-01 3.39548599E-02-1.60930874E-05    3
 2.83480628E-09 2.78195172E-14-1.40362853E+04 2.16500800E+01                   4
NC3H7O2H   8/12/15      C   3H   8O   2    0G   300.000  5000.000 1392.000    41
 1.42246236E+01 1.74340964E-02-5.97063522E-06 9.27753851E-10-5.38585168E-14    2
-2.88159737E+04-4.74357865E+01 1.35815897E+00 4.56683952E-02-2.91646368E-05    3
 9.41701313E-09-1.22337394E-12-2.41528416E+04 2.23322825E+01                   4
NC3H7O2    8/12/15      C   3H   7O   2    0G   300.000  5000.000 1390.000    31
 1.32753283E+01 1.61303126E-02-5.52348308E-06 8.58197168E-10-4.98172586E-14    2
-1.16032968E+04-4.15091215E+01 2.13311681E+00 3.96692045E-02-2.37570127E-05    3
 6.96020417E-09-7.82576856E-13-7.46687112E+03 1.92444565E+01                   4
IC3H7O2H   8/12/15      C   3H   8O   2    0G   300.000  5000.000 1405.000    41
 1.44896107E+01 1.68268026E-02-5.67601391E-06 8.72850837E-10-5.02993991E-14    2
-3.06478491E+04-5.01352281E+01 1.77384705E+00 4.75813498E-02-3.43745304E-05    3
 1.31405381E-08-2.06922904E-12-2.63458844E+04 1.77669753E+01                   4
IC3H7O2    8/12/15      C   3H   7O   2    0G   300.000  5000.000 1407.000    31
 1.35268120E+01 1.54306581E-02-5.17464218E-06 7.92548669E-10-4.55415379E-14    2
-1.33946348E+04-4.40461451E+01 2.58517502E+00 4.16107259E-02-2.92193877E-05    3
 1.08614807E-08-1.66312005E-12-9.67013161E+03 1.44731300E+01                   4
NC3H7O     8/12/15      C   3H   7O   1    0G   300.000  5000.000 1386.000    21
 1.15279177E+01 1.53775991E-02-5.23946272E-06 8.11382512E-10-4.69927603E-14    2
-9.85099867E+03-3.54233008E+01 2.57486880E+00 3.07100600E-02-1.20048836E-05    3
 3.40807108E-12 7.25275283E-13-6.20913350E+03 1.45966401E+01                   4
IC3H7O     8/12/15      C   3H   7O   1    0G   300.000  5000.000 1527.000    21
 1.19648494E+01 1.42943974E-02-4.71413211E-06 7.14027066E-10-4.07161162E-14    2
-1.17519389E+04-3.88860959E+01 2.36108410E+00 3.45650027E-02-1.94579631E-05    3
 4.71536901E-09-2.64704937E-13-8.28791395E+03 1.33112436E+01                   4
C3H6OOH1-2 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1387.000    41
 1.38088686E+01 1.43845650E-02-4.74440961E-06 7.19308280E-10-4.10654123E-14    2
-5.14352831E+03-4.20210765E+01 2.83631132E+00 3.88229894E-02-2.47944364E-05    3
 7.85644898E-09-9.58634300E-13-1.26002528E+03 1.72549973E+01                   4
C3H6OOH1-3 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1401.000    41
 1.39130757E+01 1.40218463E-02-4.55921149E-06 6.84182417E-10-3.87696213E-14    2
-3.65650518E+03-4.21532559E+01 1.74271107E+00 4.53733504E-02-3.57580373E-05    3
 1.48540053E-08-2.49981756E-12 2.32580844E+02 2.20973041E+01                   4
C3H6OOH2-1 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1393.000    41
 1.36645362E+01 1.54329764E-02-5.29285952E-06 8.23001262E-10-4.77931121E-14    2
-5.58295862E+03-4.28758364E+01 2.38465746E+00 4.42928555E-02-3.50977087E-05    3
 1.53695144E-08-2.81167824E-12-1.80979612E+03 1.69923285E+01                   4
C3H6OOH1-2O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1404.000    51
 1.91044980E+01 1.44076100E-02-4.72127814E-06 7.12631642E-10-4.05578490E-14    2
-2.50270510E+04-6.63747978E+01 3.99085043E+00 5.31865338E-02-4.28597948E-05    3
 1.77187019E-08-2.92768695E-12-2.02143526E+04 1.34150719E+01                   4
C3H6OOH1-3O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1416.000    51
 1.81661664E+01 1.47644887E-02-4.74842743E-06 7.06972467E-10-3.98305587E-14    2
-2.26256376E+04-5.93719393E+01 5.56933350E+00 4.68523421E-02-3.58917784E-05    3
 1.43314525E-08-2.29776083E-12-1.86065694E+04 7.18655005E+00                   4
C3H6OOH2-1O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1404.000    51
 1.91044980E+01 1.44076100E-02-4.72127814E-06 7.12631642E-10-4.05578490E-14    2
-2.50270510E+04-6.63747978E+01 3.99085043E+00 5.31865338E-02-4.28597948E-05    3
 1.77187019E-08-2.92768695E-12-2.02143526E+04 1.34150719E+01                   4
C3KET12   10/17/12      C   3H   6O   3    0G   300.000  5000.000 1385.000    41
 1.70187760E+01 1.32097361E-02-4.67054741E-06 7.41411770E-10-4.36869787E-14    2
-4.23572589E+04-5.92615939E+01 1.03882879E+00 5.34180080E-02-4.47684141E-05    3
 1.94651680E-08-3.45055244E-12-3.70308881E+04 2.56511209E+01                   4
C3KET13   10/17/12      C   3H   6O   3    0G   300.000  5000.000 1508.000    41
 1.73612692E+01 1.32330813E-02-4.75332110E-06 7.62529227E-10-4.52613717E-14    2
-4.06248060E+04-6.17768199E+01 4.74956819E+00 3.14080991E-02-6.83838427E-06    3
-5.67123901E-09 2.27686972E-12-3.51924570E+04 9.83753744E+00                   4
C3H51-2,3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1386.000    61
 2.12378169E+01 1.39519596E-02-4.94539222E-06 7.86381389E-10-4.63925564E-14    2
-1.92864584E+04-7.69636561E+01 2.55619708E+00 6.13504487E-02-5.23205391E-05    3
 2.28208029E-08-4.02231508E-12-1.31353414E+04 2.21043799E+01                   4
C3H52-1,3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1379.000    61
 2.02817964E+01 1.48155431E-02-5.25503386E-06 8.35963453E-10-4.93308915E-14    2
-1.80085066E+04-7.22688262E+01 4.12253742E+00 5.19553611E-02-3.83733727E-05    3
 1.45851637E-08-2.29820536E-12-1.22759164E+04 1.48367359E+01                   4
C3H5O1-2OOH-3 10/13 THERC   3H   6O   3    0G   300.000  5000.000 1432.000    31
 1.57042382E+01 1.30255692E-02-4.23544254E-06 6.35555595E-10-3.60110207E-14    2
-2.77269333E+04-5.51895464E+01-3.25001215E+00 6.65787151E-02-6.18859778E-05    3
 2.84638649E-08-5.08511634E-12-2.22371240E+04 4.30381280E+01                   4
C3H5O1-3OOH-2 10/13 THERC   3H   6O   3    0G   300.000  5000.000 1434.000    21
 1.44493479E+01 1.36372560E-02-4.25836513E-06 6.20006211E-10-3.43451580E-14    2
-2.77372360E+04-5.06099103E+01-4.43959178E+00 7.16532928E-02-7.15032351E-05    3
 3.51737842E-08-6.63682938E-12-2.27250412E+04 4.56394038E+01                   4
C3H6O1-2          A01/05C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 8.01491079E+00 1.73919953E-02-6.26027968E-06 1.01188256E-09-6.06239111E-14    2
-1.51980838E+04-1.88279964E+01 3.42806676E+00 6.25176642E-03 6.13196311E-05    3
-8.60387185E-08 3.51371393E-11-1.28446646E+04 1.04244994E+01-1.11564001E+04    4
C3H6O1-3          A11/04C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 6.80716906E+00 1.88824545E-02-6.79082475E-06 1.09713919E-09-6.57154952E-14    2
-1.36547629E+04-1.35382154E+01 5.15283752E+00-1.86401716E-02 1.29980652E-04    3
-1.58629974E-07 6.20668783E-11-1.13243512E+04 4.73561224E+00-9.75233898E+03    4
C3H6       8/12/15      C   3H   6    0    0G   298.000  6000.000 1000.000    01
 6.59032304E+00 1.52592866E-02-5.30369441E-06 8.35510888E-10-4.91215549E-14    2
-2.47481113E+02-1.15748238E+01-1.54606737E+00 4.36553128E-02-5.61392417E-05    3
 4.98421927E-08-1.84798923E-11 2.07056233E+03 2.99232495E+01                   4
C3H5-A     8/12/15      C   3H   5    0    0G   298.000  6000.000 1000.000    01
 7.37604097E+00 1.23449782E-02-4.26463882E-06 6.69045835E-10-3.92202554E-14    2
 1.77332960E+04-1.61758204E+01-3.32899442E+00 5.38423469E-02-7.65500752E-05    3
 6.35512285E-08-2.14283003E-11 2.03420628E+04 3.68038362E+01                   4
C3H5-S     8/12/15      C   3H   5    0    0G   300.000  5000.000 1390.000    11
 7.95954498E+00 1.11163183E-02-3.75197834E-06 5.77246260E-10-3.32768957E-14    2
 2.80567891E+04-1.79800372E+01 1.61793372E+00 2.44803904E-02-1.41856503E-05    3
 4.16402233E-09-4.90904795E-13 3.04291037E+04 1.66341443E+01                   4
C3H5-T     8/12/15      C   3H   5    0    0G   300.000  5000.000 1376.000    11
 7.69949212E+00 1.17803985E-02-4.07791749E-06 6.38119222E-10-3.72229675E-14    2
 2.61747145E+04-1.68305890E+01 2.29256998E+00 1.98527646E-02-6.42635654E-06    3
-5.90016395E-10 5.05491095E-13 2.85773377E+04 1.39407124E+01                   4
CC3H6                   C   3H   6O   0    0G   200.000  6000.000 1000.        1
 6.21663437E+00 1.65393591E-02-5.90075838E-06 9.48095199E-10-5.65661522E-14    2
 2.95937491E+03-1.36041009E+01 2.83278674E+00-5.21028618E-03 9.29583210E-05    3
-1.22753194E-07 4.99191366E-11 5.19520048E+03 1.08306333E+01 6.41047999E+03    4
C3H5O             KPS12 C   3H   5O   1    0G   300.000  5000.000 1402.000    01
 1.02638186E+01 1.17609932E-02-3.89837957E-06 5.92650815E-10-3.38867417E-14    2
 7.25938472E+03-2.75108651E+01 8.24068673E-01 3.46749909E-02-2.51786795E-05    3
 9.56781953E-09-1.48085302E-12 1.04203725E+04 2.28283070E+01                   4
CH2CHOCH2  8/ 8/15      C   3H   5O   1    0G   300.000  5000.000 1384.000    21
 1.20076931E+01 1.05055204E-02-3.69920541E-06 5.85629983E-10-3.44431587E-14    2
 6.97311613E+03-3.75189859E+01 1.15350351E+00 3.51253596E-02-2.50071619E-05    3
 9.00715632E-09-1.32376643E-12 1.08300872E+04 2.10606652E+01                   4
CH3CHCHO                C   3H   5O   1    0G   300.000  5000.000 1424.000    21
 1.06781476E+01 1.12805711E-02-3.89010759E-06 6.07617268E-10-3.54120848E-14    2
-7.73234209E+03-3.24971238E+01 1.47166733E+00 2.69251618E-02-1.00248013E-05    3
-1.13421435E-09 1.03416658E-12-4.04142023E+03 1.88722472E+01                   4
RALD3BG                 C   3H   5O   1     G    300.00   4000.00 1366.00      1
 .979372730E+01 .168079281E-01-.684815970E-05 .118460585E-08-.738195109E-13    2
-.875662870E+04-.294639062E+02 .667614768E+01 .261082031E-02 .280410577E-04    3
-.226802600E-07 .516442572E-11-.510504908E+04-.439698728E+01                   4
RALD3BG                 C   3H   5O   1    0G   300.000  5000.000 1424.000    21 ! CH3CHCHO
 1.06781476E+01 1.12805711E-02-3.89010759E-06 6.07617268E-10-3.54120848E-14    2
-7.73234209E+03-3.24971238E+01 1.47166733E+00 2.69251618E-02-1.00248013E-05    3
-1.13421435E-09 1.03416658E-12-4.04142023E+03 1.88722472E+01                   4
AC4H7OOH   6/17/13 THERMC   4H   8O   2    0G   300.000  5000.000 1395.000    41
 1.47661443E+01 2.12235231E-02-7.09403390E-06 1.08423759E-09-6.22145708E-14    2
-1.35617411E+04-4.77449138E+01 1.33470633E+00 5.27831440E-02-3.58861360E-05    3
 1.32495013E-08-2.06619289E-12-8.87891782E+03 2.43857336E+01                   4
C3H6OH1-2  9/ 1/12      C   3H   7O   1    0G   300.000  5000.000 1395.000    31
 1.00338281E+01 1.60227373E-02-5.41658448E-06 8.34191172E-10-4.81215988E-14    2
-1.27912397E+04-2.39034395E+01 5.05207596E-01 3.63869988E-02-2.15530901E-05    3
 6.45584786E-09-7.71267046E-13-9.26980840E+03 2.79804349E+01                   4
CH3CHCO   03/03/95 THERMC   3H   4O   1    0G   300.000  5000.000 1400.00     41
 1.00219123E+01 9.56966300E-03-3.26221644E-06 5.05231706E-10-2.92593257E-14    2
-1.42482738E+04-2.77829973E+01 1.48380119E+00 3.22203013E-02-2.70250033E-05    3
 1.20499164E-08-2.18365931E-12-1.15276540E+04 1.71552068E+01                   4
AC3H5OOH    GOLDSMITH   C   3H   6O   2    0G   298.0    6000.0   1000.000    31
 1.20838649E+01 1.47946591E-02-5.13212591E-06 8.07504999E-10-4.74394983E-14    2
-1.02184463E+04-3.36434791E+01 3.18124993E+00 4.35233041E-02-5.16277353E-05    3
 4.32011427E-08-1.57714983E-11-7.63521503E+03 1.21725683E+01                   4
C3H6OH2-1  8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1392.000    31
 1.12222277E+01 1.36444398E-02-4.51406709E-06 7.10523275E-10-4.22690392E-14    2
-1.75350136E+04-3.18911926E+01 1.09670360E+00 3.80727565E-02-2.75022497E-05    3
 1.07477493E-08-1.74895773E-12-1.40764487E+04 2.22475799E+01                   4
HOC3H6O2   9/ 1/12      C   3H   7O   3    0G   300.000  5000.000 1407.000    41
 1.56948113E+01 1.57703692E-02-5.30501726E-06 8.14307835E-10-4.68666193E-14    2
-3.24540840E+04-5.06084117E+01 2.84960487E+00 4.77244552E-02-3.60392974E-05    3
 1.43479922E-08-2.33507634E-12-2.82106103E+04 1.76478537E+01                   4
SC3H5OH    2/ 3/ 9      C   3H   6O   1    0G   300.000  5000.000 1404.000    21
 1.11222064E+01 1.27745410E-02-4.25315532E-06 6.48216484E-10-3.71190850E-14    2
-2.36690795E+04-3.41335182E+01-3.53977226E-02 4.34969453E-02-3.74479918E-05    3
 1.70906074E-08-3.13775054E-12-2.02502608E+04 2.41528201E+01                   4
IC3H5OH    8/ 1/95 THERMC   3H   6O   1    0G   300.000  5000.000 1374.00     21
 1.07381025E+01 1.31698194E-02-4.41529622E-06 6.77009837E-10-3.89608901E-14    2
-2.47298321E+04-3.13634050E+01 1.58376391E+00 3.16215366E-02-1.73664942E-05    3
 4.18927663E-09-2.79899620E-13-2.12643496E+04 1.88313766E+01                   4
C3H5OH            T06/10C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 8.72477114E+00 1.63942712E-02-5.90852993E-06 9.53262253E-10-5.70318010E-14    2
-1.90496618E+04-1.97198674E+01 3.15011905E+00 1.28538274E-02 4.28438434E-05    3
-6.67818707E-08 2.80408237E-11-1.66413668E+04 1.35066359E+01-1.48710589E+04    4
CH2CCH2OH  9/ 8/95 THERMC   3H   5O   1    0G   300.000  5000.000 1372.00     21
 9.70702027E+00 1.13972660E-02-3.77993962E-06 5.75209277E-10-3.29229125E-14    2
 9.13212884E+03-2.25012933E+01 2.88422544E+00 2.42428071E-02-1.14152268E-05    3
 1.71775334E-09 1.42177454E-13 1.17935615E+04 1.52102335E+01                   4
C3H4-P            T 2/90H  4 C  3    0    0 G   200.000  6000.00  1000.00      1
 0.60252400E+01 0.11336542E-01-0.40223391E-05 0.64376063E-09-0.38299635E-13    2
 0.19620942E+05-0.86043785E+01 0.26803869E+01 0.15799651E-01 0.25070596E-05    3
-0.13657623E-07 0.66154285E-11 0.20802374E+05 0.98769351E+01 0.22302059E+05    4
C3H4-A            L 8/89C  3 H  4    0    0 G   200.000  6000.00  1000.00      1
 0.63168722E+01 0.11133728E-01-0.39629378E-05 0.63564238E-09-0.37875540E-13    2
 0.20117495E+05-0.10995766E+02 0.26130445E+01 0.12122575E-01 0.18539880E-04    3
-0.34525149E-07 0.15335079E-10 0.21541567E+05 0.10226139E+02 0.22962267E+05    4
C3H3              T 7/11C  3 H  3    0    0 G   200.000  6000.00  1000.000     1
 7.14221719E+00 7.61902211E-03-2.67460030E-06 4.24914904E-10-2.51475443E-14    2
 3.95709594E+04-1.25848690E+01 1.35110873E+00 3.27411291E-02-4.73827407E-05    3
 3.76310220E-08-1.18541128E-11 4.07679941E+04 1.52058598E+01 4.22762135E+04    4
CC3H4             T12/81C   3H   4    0    0G   300.000  5000.00  1000.00      1
 0.66999931E+01 0.10357372E-01-0.34551167E-05 0.50652949E-09-0.26682276E-13    2
 0.30199051E+05-0.13378770E+02-0.24621047E-01 0.23197215E-01-0.18474357E-05    3
-0.15927593E-07 0.86846155E-11 0.32334137E+05 0.22729762E+02 0.3332728 E+05    4
C3H2              T12/00C  3 H  2    0    0 G   200.000  6000.00  1000.00      1
 6.67324762E+00 5.57728845E-03-1.99180164E-06 3.20289156E-10-1.91216272E-14    2
 7.57571184E+04-9.72894405E+00 2.43417332E+00 1.73013063E-02-1.18294047E-05    3
 1.02756396E-09 1.62626314E-12 7.69074892E+04 1.21012230E+01 7.83005132E+04    4
H2CCC(S)               0C   3H   2    0    0G   200.000  5000.000 1500.00    0 1
 0.64888762E+01 0.53112789E-02-0.17809490E-05 0.27252642E-09-0.15619590E-13    2
 0.63661864E+05-0.10064283E+02 0.37229726E+01 0.92589854E-02-0.23006191E-05    3
-0.10200808E-08 0.45374357E-12 0.64877289E+05 0.56865936E+01                   4
C3H2(S)                0C   3H   2    0    0G   200.000  5000.000  900.00    0 1
 0.77642570E+01 0.47112774E-02-0.16170637E-05 0.25472406E-09-0.15038572E-13    2
 0.66849672E+05-0.15098549E+02 0.52976482E+01 0.16987466E-01-0.24266517E-04    3
 0.18653681E-07-0.55763001E-11 0.67240466E+05-0.37540041E+01                   4
C3H2C                  0C   3H   2    0    0G   200.000  5000.000 1500.00    0 1
 0.65632680E+01 0.52363256E-02-0.17544830E-05 0.26866106E-09-0.15428509E-13    2
 0.56514618E+05-0.12000607E+02 0.11295888E+01 0.17287401E-01-0.11366823E-04    3
 0.34569296E-08-0.36615951E-12 0.58419080E+05 0.17331448E+02                   4
PC3H4OH-2  4/ 2/13 THERMC   3H   5O   1    0G   300.000  5000.000 1403.000    21
 1.07164095E+01 1.06066461E-02-3.51374060E-06 5.33713932E-10-3.04901511E-14    2
 4.98486803E+03-2.98329329E+01 1.42757363E+00 3.64825569E-02-3.18007132E-05    3
 1.46914605E-08-2.72331227E-12 7.80342663E+03 1.85890339E+01                   4
SC3H4OH    3/28/13      C   3H   5O   1    0G   300.000  5000.000 1407.000    21
 1.20968484E+01 9.43976596E-03-3.10773897E-06 4.69609188E-10-2.67165710E-14    2
-3.85854894E+02-3.76795997E+01 1.72870561E+00 4.41015870E-02-4.72013860E-05    3
 2.52073596E-08-5.13375710E-12 2.22720503E+03 1.43928257E+01                   4
C3H3O      2/17/14 CZHOUH   3C   3O   1     G   298.150  2000.000 1000.00      1
 4.19355696E+00 1.95625103E-02-1.22336450E-05 3.90615061E-09-5.08539231E-13    2
 3.14931737E+04 5.03216224E+00 8.75023836E-01 3.51184068E-02-3.89901356E-05    3
 2.40255750E-08-6.10883631E-12 3.20427921E+04 2.04717253E+01                   4
C3H3O2H    1/31/13      C   3H   4O   2    0G   300.000  5000.000 1385.000    31
 1.38152174E+01 8.62174763E-03-3.06710006E-06 4.88874247E-10-2.88888385E-14    2
 6.29182941E+03-4.39151257E+01 1.09787313E+00 4.22717882E-02-3.83969355E-05    3
 1.77405069E-08-3.27674312E-12 1.03592314E+04 2.30651783E+01                   4
C2HCHO     1/31/13      C   3H   2O   1    0G   300.000  5000.000 2012.000    11
 7.99952054E+00 7.07825497E-03-2.63086819E-06 4.33073185E-10-2.62003284E-14    2
 8.71863156E+03-1.57226237E+01 4.20776611E+00 1.34382727E-02-5.15442099E-06    3
-2.24570818E-11 2.74111284E-13 1.02117375E+04 5.43871873E+00                   4
C2H5CHO    8/12/15      C   3H   6O   1    0G   300.000  5000.000 1449.000    21
 1.06224453E+01 1.35569132E-02-4.60754771E-06 7.12755462E-10-4.12631683E-14    2
-2.78692266E+04-3.16628752E+01 2.18895588E+00 2.58289987E-02-6.04170058E-06    3
-3.70702654E-09 1.57131095E-12-2.42671146E+04 1.61496330E+01                   4
C2H5CO            A10/04C  3 H  5 O  1    0 G   200.000  6000.00  1000.00      1
 6.52325448E+00 1.54211952E-02-5.50898157E-06 8.85889862E-10-5.28846399E-14    2
-7.19631634E+03-5.19862218E+00 6.25722402E+00-9.17612184E-03 7.61190493E-05    3
-9.05514997E-08 3.46198215E-11-5.91616484E+03 2.23330599E+00-3.94851891E+03    4
CH2CH2CHO               C   3H   5O   1    0G   300.000  5000.000 1437.000    21
 1.00673122E+01 1.14971005E-02-3.90137798E-06 6.03029101E-10-3.48958224E-14    2
-2.75080876E+03-2.58818404E+01 2.55799036E+00 2.23391941E-02-4.89741478E-06    3
-3.58874384E-09 1.47175030E-12 4.53127696E+02 1.67016285E+01                   4
C2H3CHO           KPS12 C   3H   4O   1    0G   300.000  5000.000 1398.000    01
 9.99155394E+00 9.82348001E-03-3.31203088E-06 5.09524422E-10-2.93821890E-14    2
-1.25303509E+04-2.85168883E+01 7.33844455E-01 3.17482671E-02-2.29599468E-05    3
 8.42104232E-09-1.23613478E-12-9.38473548E+03 2.10308851E+01                   4
C2H3CO            KPS12 C   3H   3O   1    0G   300.000  5000.000 1395.000    01
 8.86032735E+00 8.48985205E-03-2.90350080E-06 4.50763986E-10-2.61524281E-14    2
 7.73489171E+03-2.06978792E+01 1.65335195E+00 2.57402596E-02-1.89009911E-05    3
 7.29174972E-09-1.16083226E-12 1.02020654E+04 1.78705872E+01                   4
CH3COCH3   8/12/15      C   3H   6O   1    0G   300.000  5000.000 1394.000    21
 8.87619308E+00 1.45700263E-02-4.84823280E-06 7.38614777E-10-4.22831194E-14    2
-3.06046242E+04-2.12730484E+01 2.20008426E+00 2.74019559E-02-1.31342003E-05    3
 2.57150371E-09-6.21509091E-14-2.79933966E+04 1.55883508E+01                   4
CH3COCH2   2/14/13 THERMC   3H   5O   1    0G   300.000  5000.000 1387.000    21
 1.09524298E+01 1.11458668E-02-3.86262877E-06 6.05088857E-10-3.53293362E-14    2
-9.60833727E+03-3.15622776E+01 1.13381826E+00 3.25095045E-02-2.10424651E-05    3
 6.64421151E-09-8.12618901E-13-6.04868361E+03 2.17158655E+01                   4
CH3COCH2O2 2/14/13 THERMC   3H   5O   3    0G   300.000  5000.000 1397.000    31
 1.65756401E+01 1.06465489E-02-3.61368681E-06 5.59053564E-10-3.23832271E-14    2
-2.42541401E+04-5.45304899E+01 1.19378141E+00 4.98027161E-02-4.17999508E-05    3
 1.74527607E-08-2.88198761E-12-1.93244224E+04 2.67877493E+01                   4
CH3COCH2O  2/ 8/13 THERMC   3H   5O   2    0G   300.000  5000.000 2002.000    21
 9.84061707E+00 1.59181106E-02-5.85164644E-06 9.56160073E-10-5.75477263E-14    2
-2.11214823E+04-2.12330791E+01 5.85960137E+00 1.78954926E-02 7.41506398E-07    3
-5.40032753E-09 1.47393197E-12-1.90714739E+04 2.70987883E+00                   4
C3KET21    2/14/13 THERMC   3H   6O   3    0G   300.000  5000.000 1394.000    41
 1.75768076E+01 1.20311704E-02-4.11633942E-06 6.40149366E-10-3.72127562E-14    2
-4.15502347E+04-6.09097100E+01-8.74352903E-01 6.12501498E-02-5.51474542E-05    3
 2.48491014E-08-4.42613472E-12-3.58060819E+04 3.59306224E+01                   4
NC4H10      8/12/15      C   4H  10    0    0G   300.000  5000.000 1392.000    31
 1.24923813E+01 2.15951935E-02-7.34277611E-06 1.13529859E-09-6.56730149E-14    2
-2.17598985E+04-4.41546866E+01-9.20862487E-02 4.69703816E-02-2.54761945E-05    3
 6.35894738E-09-5.16005946E-13-1.69556758E+04 2.49101571E+01                   4
PC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1393.000    31
 1.18547949E+01 1.96962095E-02-6.71054229E-06 1.03891144E-09-6.01513573E-14    2
 3.38182243E+03-3.72343446E+01 4.09644702E-01 4.29511341E-02-2.36582809E-05    3
 6.15744917E-09-5.64300671E-13 7.74319150E+03 2.55312526E+01                   4
SC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1682.000    31
 9.25139144E+00 2.24301385E-02-7.82648592E-06 1.23559460E-09-7.26249864E-14    2
 3.11148804E+03-2.16080436E+01 9.42662332E-01 3.77414530E-02-1.58911963E-05    3
 1.75489317E-09 2.89725750E-13 6.20542636E+03 2.42126605E+01                   4
PC4H9O                  C   4H   9O   1    0G   300.000  5000.000 1396.000    31
 1.53371588E+01 1.92789649E-02-6.56856538E-06 1.01724003E-09-5.89183466E-14    2
-1.41958782E+04-5.45071855E+01 1.84659093E+00 4.61054365E-02-2.44856516E-05    3
 5.11293268E-09-1.07538298E-13-9.09206746E+03 1.95237441E+01                   4
SC4H9O                  C   4H   9O   1    0G   300.000  5000.000 1411.000    31
 1.52130012E+01 1.90029969E-02-6.39004701E-06 9.80774402E-10-5.64493733E-14    2
-1.59888805E+04-5.43195369E+01 2.01772535E+00 4.70083969E-02-2.74726645E-05    3
 7.36290028E-09-6.30414237E-13-1.11892176E+04 1.74371746E+01                   4
PC4H9O2    8/12/15      C   4H   9O   2    0G   300.000  5000.000 1391.000    41
 1.66120049E+01 2.04752336E-02-7.01415262E-06 1.09010510E-09-6.32913959E-14    2
-1.57901735E+04-5.79272276E+01 1.80541406E+00 5.26493060E-02-3.30870383E-05    3
 1.04593484E-08-1.32305701E-12-1.03866773E+04 2.24829685E+01                   4
SC4H9O2                 C   4H   9O   2    0G   300.000  5000.000 1403.000    41
 1.68209433E+01 1.98834074E-02-6.71755569E-06 1.03411636E-09-5.96371075E-14    2
-1.75815350E+04-5.95731156E+01 2.27751066E+00 5.44334651E-02-3.82988187E-05    3
 1.42447767E-08-2.18864515E-12-1.25909100E+04 1.83237264E+01                   4
PC4H9O2H   8/12/15      C   4H  10O   2    0G   300.000  5000.000 1393.000    51
 1.75610913E+01 2.17832847E-02-7.46366287E-06 1.16012068E-09-6.73630029E-14    2
-3.30036118E+04-6.38547212E+01 1.04177717E+00 5.85996659E-02-3.84212378E-05    3
 1.28728231E-08-1.75491358E-12-2.70744200E+04 2.55179528E+01                   4
SC4H9O2H                C   4H  10O   2    0G   300.000  5000.000 1402.000    51
 1.78075939E+01 2.12546017E-02-7.20960281E-06 1.11291271E-09-6.43060022E-14    2
-3.48455718E+04-6.58011470E+01 1.44010868E+00 6.05300206E-02-4.36262678E-05    3
 1.66226146E-08-2.61556930E-12-2.92631492E+04 2.17354113E+01                   4
C4H8OOH1-2              C   4H   9O   2    0G   300.000  5000.000 1389.000    51
 1.67810269E+01 1.99677597E-02-6.85257220E-06 1.06628911E-09-6.19616154E-14    2
-9.14762760E+03-5.68667893E+01 2.91878364E+00 4.86143951E-02-2.81342168E-05    3
 7.64456491E-09-7.32889491E-13-3.94464787E+03 1.89326241E+01                   4
C4H8OOH1-3              C   4H   9O   2    0G   300.000  5000.000 1396.000    51
 1.61247782E+01 2.02420980E-02-6.88631475E-06 1.06534945E-09-6.16599545E-14    2
-9.16802012E+03-5.26575415E+01 2.46292502E+00 4.70131194E-02-2.42145198E-05    3
 4.65407810E-09 1.62198662E-14-3.95787917E+03 2.24569578E+01                   4
C4H8OOH1-4              C   4H   9O   2    0G   300.000  5000.000 1393.000    51
 1.69217927E+01 1.99305696E-02-6.85727522E-06 1.06879474E-09-6.21774931E-14    2
-7.87920857E+03-5.76630146E+01 1.35984095E+00 5.52812385E-02-3.75640846E-05    3
 1.32624209E-08-1.93623296E-12-2.34455867E+03 2.63197893E+01                   4
C4H8OOH2-1              C   4H   9O   2    0G   300.000  5000.000 1404.000    51
 1.77648250E+01 1.87777052E-02-6.36410476E-06 9.81958228E-10-5.67252066E-14    2
-9.93851667E+03-6.28169590E+01 2.32205003E+00 5.55032280E-02-3.97237996E-05    3
 1.47353739E-08-2.22481777E-12-4.67331585E+03 1.98332327E+01                   4
C4H8OOH2-3              C   4H   9O   2    0G   300.000  5000.000 1403.000    51
 1.70353922E+01 1.92729887E-02-6.50684653E-06 1.00126173E-09-5.77270961E-14    2
-1.09437234E+04-5.87403112E+01 3.30289851E+00 5.08231524E-02-3.39615358E-05    3
 1.17622237E-08-1.66012808E-12-6.13671017E+03 1.51726178E+01                   4
C4H8OOH2-4              C   4H   9O   2    0G   300.000  5000.000 1403.000    51
 1.72354039E+01 1.91946365E-02-6.49946502E-06 1.00210964E-09-5.78559962E-14    2
-9.71158144E+03-5.98986150E+01 1.82672511E+00 5.69912331E-02-4.24389492E-05    3
 1.67119278E-08-2.70635765E-12-4.54629884E+03 2.22051948E+01                   4
C4H8O1-2                C   4H   8O   1    0G   300.000  5000.000 1463.000    21
 1.41886108E+01 1.63162740E-02-5.16581368E-06 7.60173986E-10-4.24548403E-14    2
-2.02839382E+04-5.12817914E+01-4.29657099E+00 6.75906816E-02-5.89614134E-05    3
 2.59401158E-08-4.45926746E-12-1.48799944E+04 4.47755567E+01                   4
C4H8O1-3                C   4H   8O   1    0G   300.000  5000.000 1447.000    11
 1.32076917E+01 1.77467973E-02-5.69933762E-06 8.47771212E-10-4.77345874E-14    2
-2.11717546E+04-4.78386420E+01-5.37284363E+00 6.62224444E-02-5.35318273E-05    3
 2.19451842E-08-3.54479816E-12-1.54144887E+04 4.98345472E+01                   4
C4H8O1-4                C   4H   8O   1    0G   300.000  5000.000 1484.000    01
 1.22763349E+01 1.89105920E-02-6.09113637E-06 9.08066245E-10-5.12149503E-14    2
-2.92260872E+04-4.41235671E+01-7.78117916E+00 6.98405060E-02-5.45315920E-05    3
 2.13029617E-08-3.24666872E-12-2.28996340E+04 6.17620955E+01                   4
C4H8O2-3                C   4H   8O   1    0G   300.000  5000.000 1403.000    21
 1.06341771E+01 2.41442268E-02-1.13123977E-05 2.25480711E-09-1.54043041E-13    2
-2.10383343E+04-3.36763636E+01-4.48183187E+00 6.89313360E-02-6.15371646E-05    3
 2.73743747E-08-4.85890996E-12-1.68924193E+04 4.38882874E+01                   4
C4H8OOH1-2O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H8OOH1-3O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H8OOH1-4O2            C   4H   9O   4    0G   300.000  5000.000 1387.000    71
 2.26393370E+01 1.98017374E-02-6.92349554E-06 1.09100182E-09-6.39617643E-14    2
-2.75442161E+04-8.40747892E+01 2.91974455E+00 6.34948347E-02-4.29699499E-05    3
 1.42283155E-08-1.84506244E-12-2.04867301E+04 2.26279495E+01                   4
C4H8OOH2-1O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H8OOH2-3O2            C   4H   9O   4    0G   300.000  5000.000 1408.000    61
 2.19463055E+01 1.97307584E-02-6.65765380E-06 1.02424556E-09-5.90486257E-14    2
-3.07772334E+04-8.12053531E+01 3.34683971E+00 6.67468082E-02-5.25088611E-05    3
 2.14288389E-08-3.53381793E-12-2.47340662E+04 1.73189003E+01                   4
C4H8OOH2-4O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H71-2,4OOH            C   4H   9O   4    0G   300.000  5000.000 1398.000    71
 2.18629952E+01 1.99359398E-02-6.85103949E-06 1.06712096E-09-6.20561893E-14    2
-2.10042547E+04-7.80706874E+01 2.99387028E+00 6.52913914E-02-4.87958562E-05    3
 1.88107554E-08-2.95256716E-12-1.46021097E+04 2.27763716E+01                   4
C4H72-1,3OOH            C   4H   9O   4    0G   300.000  5000.000 1395.000    71
 2.14626449E+01 2.02946207E-02-6.97889021E-06 1.08750673E-09-6.32605387E-14    2
-2.22196721E+04-7.60671568E+01 3.85542428E+00 6.05523559E-02-4.18122063E-05    3
 1.46680029E-08-2.07881996E-12-1.60359412E+04 1.87734959E+01                   4
C4H72-1,4OOH            C   4H   9O   4    0G   300.000  5000.000 1387.000    71
 2.10228668E+01 2.10127561E-02-7.30349553E-06 1.14623341E-09-6.70076491E-14    2
-2.02908167E+04-7.29927491E+01 3.41714555E+00 5.89885977E-02-3.76843121E-05    3
 1.18450422E-08-1.46347291E-12-1.38437952E+04 2.27094787E+01                   4
C4H71-2,3OOH            C   4H   9O   4    0G   300.000  5000.000 1406.000    71
 2.22828679E+01 1.92253507E-02-6.52860872E-06 1.00881573E-09-5.83408336E-14    2
-2.29719991E+04-8.11231836E+01 3.30790561E+00 6.66513240E-02-5.21744859E-05    3
 2.10434152E-08-3.42495389E-12-1.67536738E+04 1.95806784E+01                   4
C4H7O1-3OOH-4           C   4H   8O   3    0G   300.000  5000.000 1418.000    31
 1.87250111E+01 1.88463312E-02-6.40165949E-06 9.89754621E-10-5.72727585E-14    2
-3.29825730E+04-7.18225468E+01-5.40949665E+00 8.05102667E-02-6.64646030E-05    3
 2.73711905E-08-4.44856733E-12-2.53005240E+04 5.56327196E+01                   4
C4H7O1-3OOH-2           C   4H   8O   3    0G   300.000  5000.000 1425.000    31
 1.97110479E+01 1.79060432E-02-6.05724664E-06 9.34110479E-10-5.39628469E-14    2
-3.52532541E+04-7.83129016E+01-4.68244067E+00 8.03419743E-02-6.67264700E-05    3
 2.74081300E-08-4.41623778E-12-2.75307409E+04 5.04193128E+01                   4
C4H7O1-2OOH-4           C   4H   8O   3    0G   300.000  5000.000 1417.000    41
 1.96187267E+01 1.77382423E-02-6.03563743E-06 9.34268374E-10-5.41073277E-14    2
-3.21917914E+04-7.50295988E+01-3.06056578E+00 7.52777235E-02-6.16382083E-05    3
 2.51520765E-08-4.05109146E-12-2.49310387E+04 4.48871201E+01                   4
C4H7O1-4OOH-2           C   4H   8O   3    0G   300.000  5000.000 1470.000    21
 1.74906412E+01 1.87794733E-02-6.05491558E-06 9.03185679E-10-5.09571870E-14    2
-4.22716632E+04-6.51860330E+01-5.17426936E+00 7.89225917E-02-6.62654132E-05    3
 2.77698767E-08-4.54377840E-12-3.53780833E+04 5.35508489E+01                   4
C4H7O1-2OOH-3           C   4H   8O   3    0G   300.000  5000.000 1435.000    41
 1.83476383E+01 1.72627711E-02-5.53440131E-06 8.21396496E-10-4.61479654E-14    2
-3.29223599E+04-6.69919656E+01-9.44964311E-01 7.31026695E-02-6.71227799E-05    3
 3.12252290E-08-5.67206759E-12-2.74510619E+04 3.25427282E+01                   4
C4H7O2-3OOH-1           C   4H   8O   3    0G   300.000  5000.000 1424.000    41
 2.03028185E+01 1.69331534E-02-5.71128715E-06 8.79005552E-10-5.07088176E-14    2
-3.43451470E+04-7.95919117E+01-3.04171082E+00 7.75254740E-02-6.55776743E-05    3
 2.74944445E-08-4.52476822E-12-2.70343494E+04 4.33136810E+01                   4
C4H72-1OOH              C   4H   8O   2    0G   300.000  5000.000 1381.000    41
 1.80122740E+01 1.70340943E-02-5.89884086E-06 9.23962123E-10-5.39539803E-14    2
-1.74585465E+04-6.55209757E+01 1.29755275E+00 5.59252255E-02-4.08890003E-05    3
 1.54880526E-08-2.42412478E-12-1.16046928E+04 2.43621382E+01                   4
NC4KET12                C   4H   8O   3    0G   300.000  5000.000 1389.000    51
 2.17577434E+01 1.64473301E-02-5.79961988E-06 9.19149624E-10-5.41037382E-14    2
-4.47115295E+04-8.37725285E+01-7.24231793E-01 7.26648886E-02-6.04779190E-05    3
 2.54348857E-08-4.30152907E-12-3.72936909E+04 3.56276963E+01                   4
NC4KET13                C   4H   8O   3    0G   300.000  5000.000 1411.000    51
 1.93085398E+01 1.73455091E-02-5.85046818E-06 9.00297947E-10-5.19274609E-14    2
-4.51023813E+04-7.04869509E+01 3.31775682E+00 5.28482064E-02-3.43211665E-05    3
 1.04562704E-08-1.12796519E-12-3.94868388E+04 1.58443308E+01                   4
NC4KET14                C   4H   8O   3    0G   300.000  5000.000 1385.000    51
 1.89231898E+01 1.82270124E-02-6.27434124E-06 9.78729382E-10-5.69844333E-14    2
-4.32508875E+04-6.78717188E+01 2.92378737E+00 5.07578011E-02-2.88360718E-05    3
 6.64649914E-09-2.83907499E-13-3.72946444E+04 1.96328202E+01                   4
NC4KET21                C   4H   8O   3    0G   300.000  5000.000 1389.000    51
 2.10786402E+01 1.61788162E-02-5.53076294E-06 8.59641186E-10-4.99535144E-14    2
-4.57563821E+04-7.88014765E+01-3.88449068E-01 6.92735051E-02-5.58731127E-05    3
 2.25791086E-08-3.63900158E-12-3.86875801E+04 3.52948090E+01                   4
NC4KET23                C   4H   8O   3    0G   300.000  5000.000 1411.000    51
 1.76877593E+01 1.84820224E-02-6.18384585E-06 9.45792334E-10-5.42981801E-14    2
-4.78594254E+04-6.06681612E+01 3.56926969E+00 5.20285891E-02-3.64134216E-05    3
 1.32007682E-08-1.93576774E-12-4.30650503E+04 1.48669401E+01                   4
NC4KET24                C   4H   8O   3    0G   300.000  5000.000 1394.000    51
 1.74146206E+01 1.92744267E-02-6.57971403E-06 1.02023879E-09-5.91418353E-14    2
-4.60663138E+04-5.80320911E+01 3.12062686E+00 5.01343936E-02-3.10194950E-05    3
 9.36512355E-09-1.07548923E-12-4.08644270E+04 1.96071994E+01                   4
C4H71-3OOH              C   4H   8O   2    0G   300.000  5000.000 1392.000    41
 1.92985494E+01 1.54534427E-02-5.25460431E-06 8.13772446E-10-4.71689947E-14    2
-1.85003480E+04-7.49926639E+01-1.50977396E+00 6.85369305E-02-5.75193633E-05    3
 2.43179107E-08-4.09788488E-12-1.18018961E+04 3.50420113E+01                   4
C4H71-3,4OOH            C   4H   9O   4    0G   300.000  5000.000 1400.000    71
 2.18394783E+01 1.98802807E-02-6.81505369E-06 1.05975117E-09-6.15560073E-14    2
-2.09468667E+04-7.79984909E+01 2.56890026E+00 6.71962184E-02-5.16999792E-05    3
 2.05770379E-08-3.32914310E-12-1.45125600E+04 2.46332539E+01                   4
C4H72-3,4OOH            C   4H   9O   4    0G   300.000  5000.000 1395.000    71
 2.14626449E+01 2.02946207E-02-6.97889021E-06 1.08750673E-09-6.32605387E-14    2
-2.22196721E+04-7.60671568E+01 3.85542428E+00 6.05523559E-02-4.18122063E-05    3
 1.46680029E-08-2.07881996E-12-1.60359412E+04 1.87734959E+01                   4
HO2CH2CHO  9/ 8/14      C   2H   4O   3    0G   300.000  5000.000 1391.000    31
 1.51554685E+01 7.57240000E-03-2.72693024E-06 4.38217189E-10-2.60434287E-14    2
-3.41419680E+04-5.01255068E+01-1.32768631E+00 5.21618601E-02-4.97327645E-05    3
 2.31272366E-08-4.20787867E-12-2.90608844E+04 3.61860491E+01                   4
IC4H10     8/12/15      C   4H  10    0    0G   300.000  5000.000 1397.000    31
 1.26422737E+01 2.14133551E-02-7.26711536E-06 1.12207226E-09-6.48434177E-14    2
-2.28293782E+04-4.66059659E+01-1.07413829E+00 5.24618320E-02-3.42407949E-05    3
 1.18817533E-08-1.73238254E-12-1.79218932E+04 2.74851665E+01                   4
IC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1397.000    31
 1.23261837E+01 1.92057770E-02-6.52063623E-06 1.00704497E-09-5.82038734E-14    2
 2.50995714E+03-4.13478742E+01 1.20802408E-01 4.73187324E-02-3.16440251E-05    3
 1.14229699E-08-1.74784642E-12 6.84032915E+03 2.44291032E+01                   4
TC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1380.000    31
 1.02682832E+01 2.09965262E-02-7.14945754E-06 1.10648358E-09-6.40498314E-14    2
 1.57542675E+02-3.00960941E+01 1.05841769E+00 3.41133739E-02-9.03156779E-06    3
-2.95313136E-09 1.41436845E-12 4.22699258E+03 2.23965051E+01                   4
TC4H9O            T08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
 1.27371509E+01 2.33707342E-02-8.50516678E-06 1.38519973E-09-8.34398061E-14    2
-1.66940150E+04-4.53156321E+01 2.77057100E+00 2.68033175E-02 4.12718360E-05    3
-7.22054739E-08 3.02642276E-11-1.27079262E+04 1.21532856E+01-1.04543262E+04    4
IC4H9O            A08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
 1.16309708E+01 2.47981574E-02-9.01550536E-06 1.46714720E-09-8.83214518E-14    2
-1.37854612E+04-3.81956151E+01 3.80297372E+00 1.56874209E-02 6.81105412E-05    3
-9.83346774E-08 3.95261902E-11-1.00832243E+04 9.78963305E+00-7.82602559E+03    4
IC4H8O     9/ 1/12      C   4H   8O   1    0G   300.000  5000.000 1394.000    21
 1.40433578E+01 2.05733637E-02-9.09519220E-06 1.73417298E-09-1.14908544E-13    2
-3.62275308E+04-6.90009668E+01-5.02573822E+00 7.51340960E-02-6.88668822E-05    3
 3.12223247E-08-5.60128818E-12-3.07481413E+04 2.96284295E+01                   4
IC3H7CHO   2/22/96 THERMC   4H   8O   1    0G   300.000  5000.000 1391.000    31
 1.37501656E+01 1.83126722E-02-6.28572629E-06 9.78250756E-10-5.68538653E-14    2
-3.26936771E+04-4.77270548E+01-2.73021382E-01 4.89696307E-02-3.12770049E-05    3
 1.00052945E-08-1.27512074E-12-2.76054737E+04 2.83451139E+01                   4
IC3H7CO    2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000    31
 1.33305736E+01 1.61873930E-02-5.56711402E-06 8.67575951E-10-5.04696549E-14    2
-1.37307001E+04-4.33958746E+01 5.03452639E-01 4.41607510E-02-2.82139091E-05    3
 8.93548675E-09-1.11327422E-12-9.07755468E+03 2.61991461E+01                   4
IC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000    31
 1.33102250E+01 1.62097959E-02-5.57575891E-06 8.69003718E-10-5.05554202E-14    2
-7.62177931E+03-4.25050854E+01 5.21481767E-01 4.43114357E-02-2.86617314E-05    3
 9.30319894E-09-1.20761563E-12-2.99677086E+03 2.68182130E+01                   4
TC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1389.000    21
 1.31013047E+01 1.66391865E-02-5.68457623E-06 8.81808351E-10-5.11290161E-14    2
-1.30638647E+04-4.42705813E+01 1.87052762E+00 4.14869677E-02-2.66815701E-05    3
 9.01531610E-09-1.27870633E-12-8.97730744E+03 1.66174178E+01                   4
IC3H5CHO                C   4H   6O   1    0G   300.000  5000.000 1396.000    21
 1.33892118E+01 1.39115420E-02-4.75820958E-06 7.38736618E-10-4.28606559E-14    2
-1.97917448E+04-4.60146004E+01 1.09372823E+00 4.43315368E-02-3.41918451E-05    3
 1.39369607E-08-2.33791460E-12-1.56745978E+04 1.94458467E+01                   4
TC3H6O2CHO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1386.00     41
 1.85534443E+01 1.68774389E-02-5.90752965E-06 9.31518085E-10-5.46345187E-14    2
-2.85447191E+04-6.82486667E+01 2.17883383E+00 5.41595832E-02-3.83435886E-05    3
 1.38308104E-08-2.04190147E-12-2.27394154E+04 2.00751264E+01                   4
IC3H5O2HCHO 8/2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00     51
 2.06288832E+01 1.48625539E-02-5.25305276E-06 8.33772951E-10-4.91277401E-14    2
-2.27589076E+04-7.82962888E+01 2.05984770E+00 5.82331716E-02-4.37672100E-05    3
 1.63249918E-08-2.43462051E-12-1.63496250E+04 2.13687921E+01                   4
TC3H6O2HCO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00     51
 2.06472678E+01 1.48526500E-02-5.25104875E-06 8.33619219E-10-4.91256069E-14    2
-2.88719869E+04-7.95951389E+01 2.03864428E+00 5.80421003E-02-4.32123528E-05    3
 1.58792094E-08-2.32209543E-12-2.24284673E+04 2.03680990E+01                   4
TC3H6OCHO  8/25/95 THERMC   4H   7O   2    0G   300.000  5000.000 1394.00     31
 1.70371287E+01 1.54400645E-02-5.28332886E-06 8.21085347E-10-4.76898429E-14    2
-2.75871941E+04-6.37271230E+01 3.70830259E-01 5.38475661E-02-3.82477565E-05    3
 1.32882237E-08-1.79228730E-12-2.18391262E+04 2.58142112E+01                   4
IC3H6CO   03/03/95 THERMC   4H   6O   1    0G   300.000  5000.000 1397.00     41
 1.32548232E+01 1.40142787E-02-4.78910215E-06 7.42924342E-10-4.30737566E-14    2
-2.00529779E+04-4.44810221E+01 2.28039055E+00 4.17016989E-02-3.25089661E-05    3
 1.37243419E-08-2.40573132E-12-1.63939712E+04 1.38187714E+01                   4
IC3H5CO                 C   4H   5O   1    0G   300.000  5000.000 1396.000    21
 1.29634401E+01 1.17954996E-02-4.04361488E-06 6.28771516E-10-3.65209867E-14    2
-8.26519462E+02-4.20562575E+01 1.87306990E+00 3.95188508E-02-3.11404053E-05    3
 1.28844447E-08-2.18165308E-12 2.85270691E+03 1.68774016E+01                   4
IC3H4CHO-A              C   4H   5O   1    0G   300.000  5000.000 1392.000    11
 1.41736959E+01 1.09161978E-02-3.69020878E-06 5.69228087E-10-3.29023246E-14    2
-1.92867979E+03-5.02663740E+01 7.64345054E-01 4.45242412E-02-3.61033720E-05    3
 1.48295287E-08-2.43809290E-12 2.44732544E+03 2.08541848E+01                   4
SC4H7OH-I         L 2/00C   4H   8O   1    0G   300.000  5000.000 1395.000    31
 1.30299481E+01 1.83782479E-02-6.18529878E-06 9.49578099E-10-5.46526348E-14    2
-3.10723026E+04-4.22891828E+01 2.70103499E+00 4.17950180E-02-2.67860575E-05    3
 9.38191037E-09-1.41171285E-12-2.73561190E+04 1.35316306E+01                   4
IC4H9O2    9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1432.000    41
 1.78793870E+01 1.82474607E-02-6.01252193E-06 9.11106794E-10-5.20018932E-14    2
-1.74569774E+04-6.61552973E+01 1.77219624E+00 5.34032789E-02-3.31041810E-05    3
 9.24465657E-09-8.01706642E-13-1.17768774E+04 2.09581481E+01                   4
TC4H9O2    9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1380.000    41
 1.80863238E+01 1.99282971E-02-6.98287309E-06 1.10171726E-09-6.46381057E-14    2
-2.04420664E+04-6.97533212E+01 2.63892371E+00 5.44717499E-02-3.75504698E-05    3
 1.40479250E-08-2.27968600E-12-1.47598933E+04 1.40325533E+01                   4
IC4H8O2H-I 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1414.000    51
 1.83915486E+01 1.73042831E-02-5.66841018E-06 8.55414265E-10-4.86781778E-14    2
-9.48569748E+03-6.67673286E+01 1.86432620E-01 6.26430177E-02-4.83690886E-05    3
 1.88657148E-08-2.91189385E-12-3.59086611E+03 2.97635367E+01                   4
IC4H8O2H-T 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1413.000    51
 1.69753885E+01 1.85198010E-02-6.09075415E-06 9.21673609E-10-5.25502501E-14    2
-1.14812757E+04-5.88259039E+01 3.84374544E+00 4.36800978E-02-2.07599526E-05    3
 2.51709167E-09 5.41306513E-13-6.50766215E+03 1.34244877E+01                   4
TC4H8O2H-I 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1379.000    51
 1.81415374E+01 1.94699499E-02-6.82750014E-06 1.07773311E-09-6.32519099E-14    2
-1.23570939E+04-6.63491602E+01 3.54378349E+00 5.25201369E-02-3.69898493E-05    3
 1.44634925E-08-2.47536050E-12-6.98183185E+03 1.27623539E+01                   4
CC4H8O     9/ 1/12      C   4H   8O   1    0G   300.000  5000.000 1431.000    11
 1.51841776E+01 1.64656666E-02-5.33483091E-06 7.98149768E-10-4.51160381E-14    2
-3.33923434E+04-7.43746988E+01-6.56746688E+00 7.87298554E-02-7.33065478E-05    3
 3.40602701E-08-6.15674656E-12-2.71582518E+04 3.80875851E+01                   4
IC4H8OOH-IO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1367.000    61
 2.24664901E+01 2.09351287E-02-7.44324128E-06 1.18589255E-09-7.00546897E-14    2
-2.94495457E+04-8.54241451E+01 4.23354857E+00 5.63088857E-02-3.15672522E-05    3
 7.79536931E-09-6.21665008E-13-2.22782534E+04 1.52623111E+01                   4
IC4H8OOH-TO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1385.000    61
 2.32464612E+01 1.88384513E-02-6.40938087E-06 9.92649459E-10-5.75275879E-14    2
-3.16533132E+04-8.88301710E+01 3.36413530E+00 6.93742776E-02-5.70416393E-05    3
 2.46040165E-08-4.32848680E-12-2.51137558E+04 1.65767339E+01                   4
TC4H8OOH-IO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1385.000    61
 2.32464612E+01 1.88384513E-02-6.40938087E-06 9.92649459E-10-5.75275879E-14    2
-3.16533132E+04-8.88301710E+01 3.36413530E+00 6.93742776E-02-5.70416393E-05    3
 2.46040165E-08-4.32848680E-12-2.51137558E+04 1.65767339E+01                   4
IC4KETII   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1387.000    51
 1.95143059E+01 1.82377395E-02-6.38908606E-06 1.00801571E-09-5.91440350E-14    2
-4.46884836E+04-7.17167584E+01 1.15501614E+00 6.10622345E-02-4.49711323E-05    3
 1.70514654E-08-2.65948602E-12-3.82747956E+04 2.69612235E+01                   4
IC4KETIT   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1388.000    51
 2.09369850E+01 1.71090955E-02-6.01892169E-06 9.52353863E-10-5.59926176E-14    2
-4.77819819E+04-8.27717611E+01 1.14243741E+00 6.33840797E-02-4.73084738E-05    3
 1.77145373E-08-2.67265475E-12-4.09366796E+04 2.34844867E+01                   4
TIC4H7Q2-I 5/ 6/96 THERMC   4H   9O   4    0G   300.000  5000.000 1400.000    71
 2.33848631E+01 1.87070035E-02-6.44021945E-06 1.00428123E-09-5.84468189E-14    2
-2.61180902E+04-8.76610135E+01 4.48426361E+00 6.61225007E-02-5.27349018E-05    3
 2.18215585E-08-3.66788946E-12-1.98906586E+04 1.26719614E+01                   4
IIC4H7Q2-I 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1394.000    71
 2.30500244E+01 1.92149194E-02-6.66622576E-06 1.04495725E-09-6.10370520E-14    2
-2.32086881E+04-8.39949885E+01 4.93055661E+00 6.05819201E-02-4.23665566E-05    3
 1.49122008E-08-2.10978665E-12-1.68415495E+04 1.36228018E+01                   4
IIC4H7Q2-T 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1377.000    71
 2.15070321E+01 2.05359839E-02-7.12383399E-06 1.11655053E-09-6.52112103E-14    2
-2.51117508E+04-7.43379783E+01 8.16274487E+00 4.34463050E-02-1.76972456E-05    3
 4.88790666E-10 9.03915465E-13-1.96501749E+04 2.62067299E-01                   4
IC4H7OOH   4/15/15      C   4H   8O   2    0G   300.000  5000.000 1386.000    41
 1.82897194E+01 1.67815784E-02-5.80668193E-06 9.08949180E-10-5.30513302E-14    2
-1.82046522E+04-6.72111342E+01 1.31851762E-01 6.19561224E-02-4.99343877E-05    3
 2.09628211E-08-3.59717924E-12-1.21399925E+04 2.93905962E+01                   4
IC4H9O2H   9/ 1/12      C   4H  10O   2    0G   300.000  5000.000 1402.000    51
 1.91651624E+01 1.93678648E-02-6.41984435E-06 9.76947752E-10-5.59299558E-14    2
-3.48790978E+04-7.42063787E+01-5.47969191E-01 6.57428787E-02-4.70123149E-05    3
 1.65991096E-08-2.27331437E-12-2.82180462E+04 3.12961385E+01                   4
TC4H9O2H   9/ 1/12      C   4H  10O   2    0G   300.000  5000.000 1382.000    51
 1.90926853E+01 2.12697804E-02-7.46252626E-06 1.17841127E-09-6.91795087E-14    2
-3.77278405E+04-7.61321196E+01 4.45573540E-01 6.66153523E-02-5.20932123E-05    3
 2.22301799E-08-4.00189859E-12-3.12260714E+04 2.37278262E+01                   4
IC4H8      8/12/15      C   4H   8    0    0G   300.000  5000.000 1392.000    21
 1.11444028E+01 1.81609265E-02-6.17791116E-06 9.55481871E-10-5.52826092E-14    2
-7.84024684E+03-3.68508829E+01 5.72478139E-02 4.17768938E-02-2.49095729E-05    3
 7.54294402E-09-9.23202212E-13-3.72166259E+03 2.35698905E+01                   4
IC4H7      8/12/15      C   4H   7    0    0G   300.000  5000.000 1384.000    11
 1.18999143E+01 1.51569859E-02-5.09995449E-06 7.83722199E-10-4.51660275E-14    2
 1.00363555E+04-4.02286635E+01-2.29578762E-01 4.17842986E-02-2.66885700E-05    3
 8.42205744E-09-1.03175361E-12 1.43946680E+04 2.54797645E+01                   4
IC4H7-I1   5/13/15      C   4H   7    0    0G   300.000  5000.000 1396.000    21
 1.11158752E+01 1.55127192E-02-5.23769366E-06 8.05998394E-10-4.64703390E-14    2
 2.19488297E+04-3.41440480E+01 9.12464579E-01 3.88654394E-02-2.57575714E-05    3
 9.07760026E-09-1.33946902E-12 2.55635553E+04 2.08634918E+01                   4
IC4H7O2           L 2/00C   4H   7O   2    0G   300.000  5000.000 1404.000    31
 1.45791608E+01 1.62136068E-02-5.26957103E-06 7.90454323E-10-4.47755051E-14    2
-1.20848042E+03-4.56459433E+01 1.43532045E+00 4.89026570E-02-3.63600970E-05    3
 1.41906420E-08-2.24557878E-12 3.09284623E+03 2.41320196E+01                   4
IC4H6OOH-I        L 2/00C   4H   7O   2    0G   300.000  5000.000 1398.000    31
 1.73601429E+01 1.42046196E-02-4.65348263E-06 7.02209785E-10-3.99552775E-14    2
-1.07509366E+03-6.12822377E+01 6.06669321E+00 3.94950065E-02-2.52721718E-05    3
 7.84485641E-09-8.98876886E-13 2.87448422E+03-3.78377026E-01                   4
CCYCCOOC-T1        THERMC   4H   7O   2    0G   300.000  5000.000 1394.000    11
 1.68269657E+01 1.64471921E-02-5.63767184E-06 8.78001611E-10-5.10959632E-14    2
-3.65710841E+03-6.74096786E+01-5.29767923E+00 6.65082201E-02-4.67054235E-05    3
 1.51029775E-08-1.74322091E-12 3.97935712E+03 5.16412476E+01                   4
C2CYCOOC-I1   7/14      C   4H   7O   2    0G   300.000  5000.000 1388.000    21
 1.89745085E+01 1.50113808E-02-5.30728309E-06 8.42454740E-10-4.96392976E-14    2
-6.93111358E+03-9.08581019E+01-2.04718031E+00 7.26608379E-02-6.82960279E-05    3
 3.27505762E-08-6.23802161E-12-3.71475599E+02 1.92056057E+01                   4
IC4H7O     4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1386.000    21
 1.33457615E+01 1.61218588E-02-5.44376403E-06 8.38199374E-10-4.83608280E-14    2
 6.11443644E+02-4.36818838E+01 1.74700687E+00 4.07783436E-02-2.44750243E-05    3
 7.06502958E-09-7.51570589E-13 4.86979233E+03 1.94535999E+01                   4
CVCYCCOC          L 2/00C   4H   6O   1    0G   300.000  5000.000 1397.000     1
 1.14363523E+01 1.63250968E-02-5.57146218E-06 8.63795613E-10-5.00701899E-14    2
-5.44653450E+03-3.87179379E+01-2.45566808E+00 4.88377067E-02-3.46186324E-05    3
 1.26590643E-08-1.88737988E-12-6.43460880E+02 3.58434061E+01                   4
CCYC2OCO          L 2/00C   4H   7O   2    0G   300.000  5000.000 1401.000    21
 1.64352871E+01 1.65843210E-02-5.71790511E-06 8.92586562E-10-5.19865043E-14    2
-1.60938498E+04-5.96946106E+01-2.97381263E+00 6.75615160E-02-5.79901709E-05    3
 2.55213006E-08-4.49991674E-12-9.93607156E+03 4.25127997E+01                   4
CCYCCOOC-I2       L 2/00C   4H   7O   2    0G   300.000  5000.000 1398.000    11
 1.63388791E+01 1.65879474E-02-5.61829108E-06 8.67331033E-10-5.01476782E-14    2
 6.66946988E+03-6.40322040E+01-4.55772603E+00 7.10221387E-02-6.05228430E-05    3
 2.61773944E-08-4.51390528E-12 1.32922215E+04 4.60828737E+01                   4
CHOIC3H6O         L 2/00C   4H   7O   2    0G   300.000  5000.000 1386.000    31
 1.55511970E+01 1.67360034E-02-5.73573457E-06 8.92095191E-10-5.18351848E-14    2
-2.50674335E+04-5.23215658E+01 2.55559437E-01 5.22086026E-02-3.72283766E-05    3
 1.36714420E-08-2.05638885E-12-1.97284649E+04 2.99210251E+01                   4
IC3H5OOCH2        L 2/00C   4H   7O   2    0G   300.000  5000.000 1410.000    41
 5.05335676E+00 3.62904388E-02-1.54012992E-05 2.74341619E-09-1.74718602E-13    2
 4.08326144E+03-2.55389509E+00-1.26548168E+00-3.61337863E-03 7.31803998E-05    3
-5.49845697E-08 1.20447492E-11 1.33108969E+04 5.33428723E+01                   4
CCYCCO-T1         L 2/00C   3H   5O   1    0G   300.000  5000.000 1389.000    11
 1.03394781E+01 1.15180335E-02-3.87496644E-06 5.95744364E-10-3.43539552E-14    2
 7.17658970E+03-2.89687593E+01-1.39311392E+00 3.81789194E-02-2.62316288E-05    3
 8.74877238E-09-1.11296763E-12 1.12534953E+04 3.41877003E+01                   4
IC4H8OH-IT              C   4H   9O   1    0G   300.000  5000.000 1391.000    41
 1.29136746E+01 2.06583409E-02-6.98445966E-06 1.07562552E-09-6.20443876E-14    2
-1.81394866E+04-3.84972088E+01 3.05275715E+00 3.93926461E-02-1.90686417E-05    3
 3.86408022E-09-1.48005244E-13-1.42263749E+04 1.60840537E+01                   4
IC4H8OH-TI              C   4H   9O   1    0G   300.000  5000.000 1402.000    41
 1.46323607E+01 1.88895981E-02-6.30561450E-06 9.62474230E-10-5.51640163E-14    2
-1.87976018E+04-4.93218793E+01 2.33169342E+00 5.13017040E-02-4.02698872E-05    3
 1.75150405E-08-3.16001727E-12-1.48318978E+04 1.55368130E+01                   4
IC4H7OH                 C   4H   8O   1    0G   300.000  5000.000 1398.000    31
 1.23304221E+01 1.83885172E-02-6.06721733E-06 9.19054723E-10-5.24036171E-14    2
-2.59452023E+04-3.67418286E+01 2.04124240E+00 4.14387207E-02-2.55228632E-05    3
 8.28133017E-09-1.10654457E-12-2.22709637E+04 1.88699473E+01                   4
IC4H8OH    2/14/95 THERMC   4H   9O   1    0G   300.000  5000.000 1376.000    41
 1.25605997E+01 2.10637488E-02-7.15019648E-06 1.10439262E-09-6.38428695E-14    2
-1.86203249E+04-3.67889430E+01 3.29612707E+00 3.47649647E-02-1.02505618E-05    3
-2.04641931E-09 1.18879408E-12-1.45627247E+04 1.58606320E+01                   4
IC4H6OH                 C   4H   7O   1    0G   300.000  5000.000 1402.000    21
 1.53490714E+01 1.38856699E-02-4.56427754E-06 6.90418690E-10-3.93540403E-14    2
-1.20164758E+04-5.55975530E+01-1.46664187E+00 6.03351671E-02-5.43112644E-05    3
 2.49299933E-08-4.52282491E-12-6.95012413E+03 3.20768458E+01                   4
TQJC4H8OH               C   4H   9O   3    0G   300.000  5000.000 1415.000    51
 2.29681617E+01 1.65162786E-02-5.50247318E-06 8.39335285E-10-4.81030625E-14    2
-4.10051460E+04-9.34897892E+01-6.43419503E-01 8.49131517E-02-8.17210578E-05    3
 3.90979927E-08-7.27092842E-12-3.42375932E+04 2.84394025E+01                   4
TQC4H8OI                C   4H   9O   3    0G   300.000  5000.000 1411.000    51
 2.13200701E+01 1.80489663E-02-6.06124072E-06 9.29740751E-10-5.34977374E-14    2
-3.12966663E+04-8.20046659E+01 7.45747835E-02 7.46499596E-02-6.42255048E-05    3
 2.80908988E-08-4.87692045E-12-2.47182737E+04 2.94511549E+01                   4
QC4H7OHP                C   4H   9O   3    0G   300.000  5000.000 1416.000    61
 2.43481084E+01 1.50316366E-02-5.01788017E-06 7.66774357E-10-4.40093220E-14    2
-3.31922320E+04-9.68211106E+01-1.27864186E+00 8.94492926E-02-8.78565423E-05    3
 4.22110919E-08-7.83450876E-12-2.58975226E+04 3.53963909E+01                   4
TQC4H7OHI         L 2/00C   4H   9O   3    0G   300.000  5000.000 1404.000    61
 2.08281225E+01 1.81675094E-02-6.12943202E-06 9.43194119E-10-5.43937008E-14    2
-3.37386684E+04-7.74823720E+01 2.55843807E+00 6.37086077E-02-4.97169945E-05    3
 1.99225109E-08-3.21373436E-12-2.77526909E+04 1.95001368E+01                   4
CCY(CCO)COH             C   4H   8O   2    0G   300.000  5000.000 1412.000    31
 1.91884885E+01 1.56255714E-02-5.22569800E-06 7.99171074E-10-4.58832445E-14    2
-4.71120302E+04-7.84579023E+01-7.10048774E+00 9.53371808E-02-9.78701612E-05    3
 4.90005646E-08-9.41685766E-12-3.98987202E+04 5.60924667E+01                   4
C2CY(COC)OH             C   4H   8O   2    0G   300.000  5000.000 1393.000    31
 1.56829970E+01 1.92910506E-02-6.63718495E-06 1.03441014E-09-6.01715267E-14    2
-4.10598236E+04-5.85686221E+01 5.92324183E-01 5.52429007E-02-4.02419018E-05    3
 1.57152217E-08-2.57388393E-12-3.58241476E+04 2.23378086E+01                   4
IQJC4H8OH         L 2/00C   4H   9O   3    0G   300.000  5000.000 1410.000    51
 2.11752212E+01 1.75144254E-02-5.73227292E-06 8.63386596E-10-4.90282414E-14    2
-3.98881576E+04-8.19187015E+01 1.81448831E+00 7.47452750E-02-7.10895172E-05    3
 3.44973679E-08-6.54646593E-12-3.44023586E+04 1.77380434E+01                   4
IC3H6OHCHO              C   4H   8O   2    0G   300.000  5000.000 1393.000    41
 1.60254376E+01 1.85402212E-02-6.36973877E-06 9.91732739E-10-5.76472640E-14    2
-5.50198923E+04-5.83074874E+01 1.84080874E+00 5.29601347E-02-3.94261774E-05    3
 1.59063430E-08-2.69565279E-12-5.01437169E+04 1.75482756E+01                   4
IQC4H8OT                C   4H   9O   3    0G   300.000  5000.000 1405.000    51
 2.04823628E+01 1.82966721E-02-6.04413378E-06 9.16380548E-10-5.22866551E-14    2
-2.94287153E+04-7.53563247E+01 3.72211529E+00 6.42864861E-02-5.52809053E-05    3
 2.50036630E-08-4.53471908E-12-2.43110525E+04 1.21981167E+01                   4
IQC4H7OHT               C   4H   9O   3    0G   300.000  5000.000 1413.000    61
 2.19945886E+01 1.62011186E-02-5.23758492E-06 7.81898296E-10-4.41125515E-14    2
-3.07383725E+04-8.16613568E+01 3.58900054E+00 7.25591129E-02-7.14080484E-05    3
 3.55250907E-08-6.84991795E-12-2.57241250E+04 1.23766657E+01                   4
CCY(CCOC)OH       L 2/00C   4H   8O   2    0G   300.000  5000.000 1404.000    21
 1.43404718E+01 1.98311504E-02-6.60657660E-06 1.00779570E-09-5.77614335E-14    2
-4.30959414E+04-5.30535015E+01-2.84914896E+00 6.23736856E-02-4.70326536E-05    3
 1.84908286E-08-2.94976027E-12-3.74257004E+04 3.83163588E+01                   4
CH2COHCH2OOH            C   3H   6O   3    0G   300.000  5000.000 1398.000    41
 1.87971268E+01 1.12783442E-02-3.90789058E-06 6.12064651E-10-3.57305453E-14    2
-3.61154867E+04-6.94914300E+01-3.89823383E-01 7.01531131E-02-7.42036788E-05    3
 3.84181056E-08-7.63555985E-12-3.07879938E+04 2.86873505E+01                   4
TC3H6OH    8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1392.000    31
 1.12222277E+01 1.36444398E-02-4.51406709E-06 7.10523275E-10-4.22690392E-14    2
-1.75350136E+04-3.18911926E+01 1.09670360E+00 3.80727565E-02-2.75022497E-05    3
 1.07477493E-08-1.74895773E-12-1.40764487E+04 2.22475799E+01                   4
TQC4H7OHIO2             C   4H   9O   5    0G   300.000  5000.000 1402.000    71
 2.82564819E+01 1.66969871E-02-5.67314614E-06 8.78350442E-10-5.09090253E-14    2
-5.66017464E+04-1.15147927E+02 3.17336206E+00 7.94005900E-02-6.51165712E-05    3
 2.62035931E-08-4.13406290E-12-4.84943162E+04 1.77867184E+01                   4
TQC4H7OHTO2             C   4H   9O   5    0G   300.000  5000.000 1402.000    71
 2.82564819E+01 1.66969871E-02-5.67314614E-06 8.78350442E-10-5.09090253E-14    2
-5.66017464E+04-1.15147927E+02 3.17336206E+00 7.94005900E-02-6.51165712E-05    3
 2.62035931E-08-4.13406290E-12-4.84943162E+04 1.77867184E+01                   4
TQC4H7OHIQ-I            C   4H   9O   5    0G   300.000  5000.000 1384.000    71
 2.88466964E+01 1.66289773E-02-5.74301906E-06 8.98791324E-10-5.24794891E-14    2
-4.69249234E+04-1.19117836E+02 6.09881562E+00 6.93745451E-02-5.12049498E-05    3
 1.81276221E-08-2.46329781E-12-3.91393707E+04 2.93862639E+00                   4
TQC4H7OHIQ-P            C   4H   9O   5    0G   300.000  5000.000 1400.000    81
 2.81439191E+01 1.63524649E-02-5.54998081E-06 8.58603978E-10-4.97359401E-14    2
-4.84502814E+04-1.11572783E+02 3.36947511E+00 7.96855226E-02-6.74365765E-05    3
 2.82233283E-08-4.65270820E-12-4.05567534E+04 1.92726029E+01                   4
IC3H5COHQ               C   4H   8O   3    0G   300.000  5000.000 1504.000    51
 2.07387831E+01 1.58360934E-02-5.27614462E-06 8.05932218E-10-4.62682425E-14    2
-4.41821241E+04-7.94239893E+01 2.64360992E+00 5.72485066E-02-3.95907807E-05    3
 1.27775635E-08-1.47241476E-12-3.80099993E+04 1.77322273E+01                   4
CH2CQCOHQ  7/ 1/14      C   3H   6O   5    0G   300.000  5000.000 1418.000    61
 3.86574091E+01 4.83815026E-04-2.10413843E-07 3.81490832E-11-2.46187754E-15    2
-6.56392184E+04-1.61083579E+02-1.61171759E+01 1.78866440E-01-2.16751308E-04    3
 1.15450289E-07-2.27163078E-11-5.21165145E+04 1.14441286E+02                   4
IC3H5Q                  C   3H   6O   2    0G   300.000  5000.000 1397.000    31
 1.43424294E+01 1.28053632E-02-4.40584813E-06 6.86848148E-10-3.99675209E-14    2
-1.65261025E+04-4.89934539E+01 1.32903007E+00 4.49170722E-02-3.51235127E-05    3
 1.41982181E-08-2.33335008E-12-1.21898396E+04 2.02696565E+01                   4
CH3COCHO                C   3H   4O   2    0G   300.000  5000.000 1381.000    21
 1.14371190E+01 1.06773624E-02-3.68967757E-06 5.77006752E-10-3.36532201E-14    2
-3.78079398E+04-3.25054087E+01 2.08731049E+00 3.09032484E-02-1.98794164E-05    3
 6.26174519E-09-7.69945504E-13-3.43989451E+04 1.82839639E+01                   4
IC3H5OCH2  6/ 2/14 CZHOUH   7C   4O   1     G   298.150  2000.000 1000.00      1
 6.64731727E+00 3.08190709E-02-1.73209320E-05 5.01099629E-09-6.00089387E-13    2
 1.70679921E+03-5.91214819E+00-2.14798958E+00 7.00225553E-02-8.21595440E-05    3
 5.22589946E-08-1.34176532E-11 3.26474773E+03 3.55145589E+01                   4
IC4H7OOCH3              C   5H  10O   2    0G   300.000  5000.000 1386.000    51
 1.95896715E+01 2.31057369E-02-8.02911330E-06 1.25969946E-09-7.36169360E-14    2
-1.80069088E+04-7.34192482E+01 1.26784161E+00 6.82442475E-02-5.30807931E-05    3
 2.27496198E-08-4.11475065E-12-1.16767937E+04 2.44900544E+01                   4
IC4H7OOIC4H7            C   8H  14O   2    0G   300.000  5000.000 1390.000    71
 2.80447245E+01 3.27505220E-02-1.13220177E-05 1.77027767E-09-1.03211988E-13    2
-1.72683337E+04-1.15134796E+02-2.07881710E-01 1.04075647E-01-8.33973077E-05    3
 3.60897624E-08-6.47906520E-12-7.79062693E+03 3.50446555E+01                   4
C4H8-1                  C   4H   8    0    0G   300.000  5000.000 1388.000    21
 1.10189295E+01 1.82714177E-02-6.21801907E-06 9.62038611E-10-5.56791341E-14    2
-5.80998818E+03-3.47942287E+01 1.62599556E-01 4.01052746E-02-2.18038592E-05    3
 5.47070727E-09-4.54073315E-13-1.65402601E+03 2.48169258E+01                   4
C4H8-2     8/12/15      C   4H   8    0    0G   300.000  5000.000 1383.000    21
 1.08652083E+01 1.84123129E-02-6.26886673E-06 9.70205962E-10-5.61638967E-14    2
-7.09625867E+03-3.51547481E+01 1.30795510E+00 3.53136624E-02-1.51866126E-05    3
 1.64112363E-09 3.44257620E-13-3.19767852E+03 1.81594717E+01                   4
C4H71-1                 C   4H   7    0    0G   300.000  5000.000 1390.000    21
 1.10531750E+01 1.55668782E-02-5.25853044E-06 8.09627095E-10-4.67015477E-14    2
 2.39455759E+04-3.31548457E+01 8.97231085E-01 3.77003788E-02-2.33194855E-05    3
 7.38468124E-09-9.50027900E-13 2.76498158E+04 2.19835413E+01                   4
C4H71-2                 C   4H   7    0    0G   300.000  5000.000 1381.000    21
 1.07105686E+01 1.63539126E-02-5.63688038E-06 8.79591989E-10-5.12098725E-14    2
 2.21011255E+04-3.15300308E+01 1.56405993E+00 3.32162309E-02-1.59178310E-05    3
 2.92637814E-09-3.02645386E-14 2.57966120E+04 1.93052496E+01                   4
C4H71-3    1/13/16      C   4H   7    0    0G   300.000  5000.000 1367.000    11
 1.16977564E+01 1.53404517E-02-5.16928607E-06 7.95431212E-10-4.58914150E-14    2
 1.07395001E+04-3.82992966E+01 9.40350126E-01 3.56830321E-02-1.74384567E-05    3
 2.78964567E-09 1.78068599E-13 1.49303203E+04 2.11349333E+01                   4
C4H71-4                 C   4H   7    0    0G   300.000  5000.000 1389.000    21
 1.03875084E+01 1.63677264E-02-5.58416036E-06 8.65388736E-10-5.01415385E-14    2
 1.93282846E+04-2.86081068E+01 5.36903096E-01 3.66356251E-02-2.07814610E-05    3
 5.74895154E-09-6.05742821E-13 2.30645349E+04 2.53369983E+01                   4
C4H72-2    8/12/15      C   4H   7    0    0G   300.000  5000.000 1378.000    21
 1.05359634E+01 1.65535631E-02-5.71669066E-06 8.93155269E-10-5.20432637E-14    2
 2.08161211E+04-3.11046229E+01 2.46499885E+00 2.94957335E-02-1.08904521E-05    3
 9.17747264E-11 5.46417906E-13 2.42904093E+04 1.44728237E+01                   4
C4H71-O    4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1395.000    21
 1.53137780E+01 1.43427017E-02-4.81625517E-06 7.39574839E-10-4.26140814E-14    2
-7.29342884E+02-5.52937859E+01-1.60619192E+00 5.58562682E-02-4.35595767E-05    3
 1.70589279E-08-2.65635180E-12 4.85090326E+03 3.47112559E+01                   4
PC4H8OH-2               C   4H   9O   1    0G   300.000  5000.000 1396.000    41
 1.47198620E+01 1.93691825E-02-6.59356634E-06 1.02018538E-09-5.90410746E-14    2
-1.53023402E+04-4.85296396E+01 1.89476538E+00 4.87803114E-02-3.26702980E-05    3
 1.17119949E-08-1.77100238E-12-1.07455371E+04 2.06226225E+01                   4
SC4H8OH-1               C   4H   9O   1    0G   300.000  5000.000 1405.000    41
 1.50517242E+01 1.84748629E-02-6.15327969E-06 9.38017339E-10-5.37214281E-14    2
-1.71974443E+04-5.03733848E+01 1.78282749E+00 5.18872497E-02-3.89600849E-05    3
 1.57818686E-08-2.64133852E-12-1.28305019E+04 2.00308244E+01                   4
SC4H8OH-3               C   4H   9O   1    0G   300.000  5000.000 1403.000    41
 1.42453780E+01 1.89491000E-02-6.27403528E-06 9.52692609E-10-5.44157896E-14    2
-1.81803642E+04-4.56206494E+01 1.93185505E+00 4.79506224E-02-3.23719194E-05    3
 1.16232751E-08-1.72498918E-12-1.39431370E+04 2.03995003E+01                   4
C4H71-3OH               C   4H   8O   1    0G   300.000  5000.000 1385.000    31
 1.42401634E+01 1.83038695E-02-6.37213444E-06 1.00099740E-09-5.85511411E-14    2
-2.68183960E+04-4.83949774E+01 7.16707858E-02 5.04772909E-02-3.50356983E-05    3
 1.30539199E-08-2.07783174E-12-2.16983717E+04 2.82072724E+01                   4
C4H71-4OH               C   4H   8O   1    0G   300.000  5000.000 1396.000    31
 1.33437331E+01 1.82063693E-02-6.15150719E-06 9.47318576E-10-5.46543216E-14    2
-2.48479001E+04-4.27998774E+01-2.12276307E-01 4.86358034E-02-3.17241965E-05    3
 1.04986646E-08-1.39007078E-12-2.00365173E+04 3.04092052E+01                   4
C4H71-1OH               C   4H   8O   1    0G   300.000  5000.000 1402.000    31
 1.42586569E+01 1.71932504E-02-5.74956414E-06 8.79089774E-10-5.04586493E-14    2
-2.78051048E+04-4.96581579E+01-4.65981165E-01 5.56573217E-02-4.50578305E-05    3
 1.93726056E-08-3.38967639E-12-2.31007894E+04 2.79744544E+01                   4
C4H71-2OH               C   4H   8O   1    0G   300.000  5000.000 1404.000    31
 1.50658194E+01 1.65276030E-02-5.52197706E-06 8.43591643E-10-4.83870716E-14    2
-2.99737946E+04-5.53405024E+01-1.28560619E+00 6.35758020E-02-5.85328191E-05    3
 2.80452715E-08-5.32187122E-12-2.51538600E+04 2.93802791E+01                   4
C4H72-1OH               C   4H   8O   1    0G   300.000  5000.000 1367.000    31
 1.32893235E+01 1.93843938E-02-6.80733358E-06 1.07559847E-09-6.31698641E-14    2
-2.58627911E+04-4.34782359E+01 2.94637661E+00 3.45852975E-02-1.10024787E-05    3
-1.33281467E-09 9.54964043E-13-2.12241816E+04 1.55037145E+01                   4
C4H72-2OH               C   4H   8O   1    0G   300.000  5000.000 1402.000    31
 1.49411596E+01 1.66289929E-02-5.55627511E-06 8.48898851E-10-4.86949390E-14    2
-3.12496851E+04-5.51730870E+01-1.84033728E-01 5.90104774E-02-5.22507028E-05    3
 2.44135801E-08-4.56518659E-12-2.66717960E+04 2.36075268E+01                   4
SQC4H8OP                C   4H   9O   3    0G   300.000  5000.000 1421.000    51
 2.02482113E+01 1.90403096E-02-6.41818812E-06 9.86791658E-10-5.68666168E-14    2
-2.70686177E+04-7.43734665E+01 3.92966105E+00 5.67740736E-02-3.88077818E-05    3
 1.31554059E-08-1.72822772E-12-2.14649445E+04 1.32313419E+01                   4
PQC4H8OS                C   4H   9O   3    0G   300.000  5000.000 1403.000    51
 1.99993833E+01 1.96391125E-02-6.70755815E-06 1.04036085E-09-6.03187960E-14    2
-2.71257575E+04-7.31284601E+01 2.68979886E+00 6.10664073E-02-4.46910607E-05    3
 1.68939056E-08-2.59692346E-12-2.12460925E+04 1.94271757E+01                   4
PQC4H7OHS-3             C   4H   9O   3    0G   300.000  5000.000 1404.000    61
 1.89703648E+01 1.96512375E-02-6.61522830E-06 1.01590849E-09-5.84889733E-14    2
-2.92876345E+04-6.40682635E+01 3.14058820E+00 5.94343278E-02-4.55414505E-05    3
 1.85507067E-08-3.10109441E-12-2.40765022E+04 1.99412365E+01                   4
NC4KET12OH              C   4H   8O   2    0G   300.000  5000.000 1384.000    41
 1.68650782E+01 1.83319076E-02-6.41389893E-06 1.01105283E-09-5.92858731E-14    2
-5.27353126E+04-5.97188408E+01 5.20269850E-01 5.40316915E-02-3.57074151E-05    3
 1.18022134E-08-1.57485744E-12-4.67781081E+04 2.89999061E+01                   4
SQC4H7OHS-4             C   4H   9O   3    0G   300.000  5000.000 1414.000    61
 2.06664415E+01 1.78772156E-02-5.93193686E-06 9.02005813E-10-5.15691990E-14    2
-3.04132233E+04-7.44595459E+01 3.37952725E+00 6.50949152E-02-5.59109752E-05    3
 2.49644089E-08-4.44896795E-12-2.51501593E+04 1.58596901E+01                   4
SQC4H8OS                C   4H   9O   3    0G   300.000  5000.000 1424.000    51
 2.05363895E+01 1.85261859E-02-6.18257770E-06 9.44045247E-10-5.41390400E-14    2
-2.90453556E+04-7.66224497E+01 3.45579406E+00 6.10420456E-02-4.64106547E-05    3
 1.80687264E-08-2.81124474E-12-2.34835698E+04 1.39991890E+01                   4
NC4KET23OH    7/27/15   C   4H   8O   2    0G   300.000  5000.000 1386.000    41
 1.54636087E+01 1.92120108E-02-6.64681122E-06 1.03988604E-09-6.06552757E-14    2
-5.57292725E+04-5.19147488E+01 1.64761234E+00 4.74122084E-02-2.72508571E-05    3
 7.25755846E-09-6.68682869E-13-5.04946247E+04 2.37800424E+01                   4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
 1.12685690E+01 2.01724820E-02-7.41925667E-06 1.21275519E-09-7.30115348E-14    2
 2.13876442E+03-3.15208064E+01 5.16434924E+00 2.53427725E-02-1.39669041E-06    3
-6.00713944E-09 1.76696879E-12 5.03210693E+03 4.37441148E+00                   4
C4H6-1            L10/93C  4.H  6.   0.   0.G   200.000  6000.000 1000.        1
 7.81179394E+00 1.79733772E-02-6.61044149E-06 1.05501491E-09-6.19297169E-14    2
 1.61770171E+04-1.59658015E+01 2.42819263E+00 2.49821955E-02 6.27370548E-06    3
-2.61747866E-08 1.26585079E-11 1.80248564E+04 1.36683982E+01 1.98688798E+04    4
AC3H5OCH2  9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1397.000    31
 1.19880368E+01 1.70263516E-02-5.78617265E-06 8.94150465E-10-5.16994613E-14    2
 3.48367473E+03-3.35860630E+01 1.20089076E+00 4.24760987E-02-2.94114641E-05    3
 1.11824860E-08-1.81309530E-12 7.26792055E+03 2.43628654E+01                   4
C5H10-2    9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1385.000    31
 1.39425521E+01 2.28734997E-02-7.77800113E-06 1.20284861E-09-6.95972140E-14    2
-1.12165700E+04-4.95379542E+01 5.90528835E-01 4.85275113E-02-2.43231598E-05    3
 4.86096027E-09-1.13099201E-13-5.99777644E+03 2.41816377E+01                   4
CC5H10     9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1394.000    31
 1.44242929E+01 2.26454984E-02-7.73646334E-06 1.19999861E-09-6.95711276E-14    2
-1.14981027E+04-5.30391197E+01-9.64397004E-01 5.68482691E-02-3.66324275E-05    3
 1.23008921E-08-1.71392531E-12-5.93502026E+03 3.02998433E+01                   4
C6H10D24                C   6H  10    0    0G   300.000  5000.000 1393.000    31
 1.67662657E+01 2.32109616E-02-7.93355119E-06 1.23101995E-09-7.13892514E-14    2
-2.93324539E+03-6.44104411E+01-3.63783422E-01 6.36719104E-02-4.53090160E-05    3
 1.73368393E-08-2.79133016E-12 3.04087286E+03 2.75469470E+01                   4
C5H91-3    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1390.000    21
 1.39593933E+01 2.09180210E-02-7.14307074E-06 1.10781333E-09-6.42268160E-14    2
 7.02651017E+03-5.03103610E+01-4.68159636E-01 5.13472600E-02-3.05648794E-05    3
 8.82809744E-09-9.61458255E-13 1.23781446E+04 2.83587835E+01                   4
C5H92-4    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1384.000    21
 1.35637956E+01 2.11621316E-02-7.20826071E-06 1.11611006E-09-6.46370085E-14    2
 5.82258629E+03-4.87323606E+01 2.55028348E-01 4.69860501E-02-2.40447582E-05    3
 4.89006694E-09-1.15557679E-13 1.09775103E+04 2.46226810E+01                   4
C5H92-5    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1386.000    31
 1.32988753E+01 2.09845923E-02-7.14999241E-06 1.10717347E-09-6.41183619E-14    2
 1.39270369E+04-4.32758927E+01 9.96363945E-01 4.49148898E-02-2.30951498E-05    3
 5.01698735E-09-2.38646470E-13 1.87161506E+04 2.45616052E+01                   4
C5H91-4    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1387.000    31
 1.29229725E+01 2.10931621E-02-7.14227112E-06 1.10137556E-09-6.35983966E-14    2
 1.38192408E+04-4.00293126E+01 1.58797615E+00 4.01577239E-02-1.50062687E-05    3
-3.94608061E-10 1.02064182E-12 1.84683983E+04 2.34273438E+01                   4
C5H91-5    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1391.000    31
 1.37334869E+01 2.07003006E-02-7.06962737E-06 1.09638953E-09-6.35591113E-14    2
 1.51176253E+04-4.50794850E+01 2.07676634E-01 4.96049077E-02-3.00621602E-05    3
 9.19962077E-09-1.13246061E-12 2.01251866E+04 2.85856261E+01                   4
C5H9O2-4   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1376.000    31
 1.73707371E+01 2.09044827E-02-7.30723872E-06 1.15106814E-09-6.74601377E-14    2
-5.48020434E+03-6.50109045E+01 3.38899911E+00 4.71704753E-02-2.40389823E-05    3
 4.99166621E-09-2.03242522E-13 1.15232772E+02 1.25183625E+01                   4
SC3H5OCH2-1             C   4H   7O   1    0G   300.000  5000.000 1382.000    31
 1.47022035E+01 1.55342107E-02-5.45701052E-06 8.62544885E-10-5.06734446E-14    2
 1.81294800E+03-5.05120353E+01 2.35694446E-01 4.67367652E-02-3.04880689E-05    3
 9.75216148E-09-1.23281228E-12 7.11668364E+03 2.81378517E+01                   4
NC4KET21OH              C   4H   8O   2    0G   300.000  5000.000 1507.000    41
 1.52252911E+01 1.86615017E-02-6.30658772E-06 9.72355897E-10-5.61770184E-14    2
-5.34759661E+04-5.00397269E+01 5.46677192E+00 3.01119974E-02-2.59548850E-06    3
-7.61700554E-09 2.55573161E-12-4.89909104E+04 6.33307684E+00                   4
C2H5CHOHCO              C   4H   7O   2    0G   300.000  5000.000 1389.000    41
 1.82917246E+01 1.48007410E-02-5.24974573E-06 8.35220286E-10-4.92942253E-14    2
-3.36703722E+04-7.12363783E+01-2.44749259E+00 6.46308488E-02-5.10457937E-05    3
 1.99850773E-08-3.12214490E-12-2.66670442E+04 3.95566556E+01                   4
CH3COCOHCH3             C   4H   7O   2    0G   300.000  5000.000 1395.000    41
 1.65624631E+01 1.59037217E-02-5.54554278E-06 8.72274939E-10-5.10735025E-14    2
-3.65884887E+04-6.10833920E+01-1.65607674E+00 6.08409982E-02-4.85215440E-05    3
 1.97794382E-08-3.26305133E-12-3.05158227E+04 3.58911868E+01                   4
C2H4COCH2OH             C   4H   7O   2    0G   300.000  5000.000 1462.000    41
 1.40828195E+01 1.76833414E-02-6.09759192E-06 9.52794521E-10-5.55571628E-14    2
-3.37518398E+04-4.08944306E+01 7.98874348E+00 1.41152447E-02 1.86299924E-05    3
-1.99223089E-08 5.12983835E-12-2.98706372E+04-1.87192030E+00                   4
CH3COHCO   9/24/15      C   3H   4O   2    0G   300.000  5000.000 1410.000    21
 1.50110709E+01 7.26697312E-03-2.42872486E-06 3.71246886E-10-2.13068531E-14    2
-3.87354954E+04-5.41005540E+01 8.25855205E-01 5.22217422E-02-5.66992291E-05    3
 2.94815948E-08-5.81714952E-12-3.50157127E+04 1.78488731E+01                   4
CH2COHCHO  9/24/15      C   3H   4O   2    0G   300.000  5000.000 1406.000    21
 1.40200417E+01 7.95092924E-03-2.63244516E-06 3.99896432E-10-2.28538120E-14    2
-3.76808145E+04-4.80457990E+01 5.76639663E-02 5.16589617E-02-5.49773816E-05    3
 2.83487148E-08-5.57464421E-12-3.39594513E+04 2.29757289E+01                   4
NC4KET13OH-2            C   4H   8O   4    0G   300.000  5000.000 1395.000    61
 2.25434165E+01 1.76377030E-02-6.14926113E-06 9.67201484E-10-5.66321794E-14    2
-6.59724022E+04-8.48522697E+01 2.13332105E+00 6.69840817E-02-5.19672275E-05    3
 2.03864253E-08-3.22074763E-12-5.90962942E+04 2.40964870E+01                   4
NC4KET24OH-1            C   4H   8O   4    0G   300.000  5000.000 1672.000    61
 1.76639507E+01 2.38921914E-02-8.87612081E-06 1.46065294E-09-8.83476797E-14    2
-6.36561283E+04-5.60405234E+01 7.17383002E+00 3.72830917E-02-7.30000099E-06    3
-5.42423663E-09 1.94298976E-12-5.91469605E+04 3.98040888E+00                   4
NC4KET24OH-3            C   4H   8O   4    0G   300.000  5000.000 1392.000    61
 2.02237496E+01 1.94540798E-02-6.73928381E-06 1.05529414E-09-6.15931037E-14    2
-6.68651215E+04-6.99676945E+01 2.60979522E+00 6.11530456E-02-4.50409252E-05    3
 1.73313054E-08-2.75573967E-12-6.07708447E+04 2.44892030E+01                   4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
 2.15163584E+01 1.55811846E-02-5.27569793E-06 8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00 7.72727339E-02-6.79667571E-05    3
 2.98158102E-08-5.16343458E-12-3.01649655E+04 4.06810164E+01                   4
C4H6OHOOH2-2-1          C   4H   8O   3    0G   300.000  5000.000 1396.000    51
 2.16656460E+01 1.59965487E-02-5.52214578E-06 8.62740322E-10-5.02768063E-14    2
-4.14875437E+04-8.39377540E+01 4.72576793E-02 7.85787048E-02-7.68006410E-05    3
 3.79206120E-08-7.33203833E-12-3.51140091E+04 2.80064858E+01                   4
C4H6OHOOH1-3-4          C   4H   8O   3    0G   300.000  5000.000 1391.000    51
 1.93445152E+01 1.82185729E-02-6.34491630E-06 9.97097673E-10-5.83420009E-14    2
-3.79952136E+04-6.88144861E+01 9.44277749E-01 6.34330602E-02-4.99455695E-05    3
 2.05720571E-08-3.48143957E-12-3.17827282E+04 2.92923796E+01                   4
C4H6OHOOH1-2-3          C   4H   8O   3    0G   300.000  5000.000 1403.000    51
 2.32793098E+01 1.38280934E-02-4.61330737E-06 7.05319574E-10-4.05174739E-14    2
-4.26348237E+04-9.51979841E+01-2.88475927E+00 9.16099207E-02-9.37152074E-05    3
 4.66406895E-08-8.92736049E-12-3.52899912E+04 3.92851633E+01                   4
HOCH2CHO   9/24/15      C   2H   4O   2    0G   300.000  5000.000 1680.000    21
 7.99598542E+00 1.20664034E-02-4.43693399E-06 7.25167046E-10-4.36535460E-14    2
-4.09020567E+04-1.33754312E+01 4.35084369E+00 1.50412895E-02-5.95083030E-07    3
-3.75736217E-09 1.09353598E-12-3.91654526E+04 8.09610238E+00                   4
C4H71-4OOH              C   4H   8O   2    0G   300.000  5000.000 1392.000    41
 1.59871304E+01 1.86028119E-02-6.40003189E-06 9.97531711E-10-5.80334203E-14    2
-1.70152141E+04-5.46227137E+01 1.31653247E+00 5.16546159E-02-3.47310922E-05    3
 1.20405755E-08-1.71650639E-12-1.17754576E+04 2.46384545E+01                   4
C4H71-4O2  9/25/15      C   4H   7O   2    0G   300.000  5000.000 1390.000    31
 1.50240251E+01 1.72860962E-02-5.94297061E-06 9.25861430E-10-5.38461748E-14    2
 1.92460667E+02-4.85941022E+01 2.09042625E+00 4.57130080E-02-2.94815830E-05    3
 9.69604853E-09-1.30061388E-12 4.88932667E+03 2.15456077E+01                   4
C4H61-3OOH4             C   4H   7O   2    0G   300.000  5000.000 1391.000    31
 1.55818475E+01 1.69176098E-02-5.84009100E-06 9.12401042E-10-5.31699330E-14    2
 1.20753065E+01-5.36683745E+01 1.00320366E+00 4.99893791E-02-3.43100656E-05    3
 1.20104294E-08-1.71132691E-12 5.17744264E+03 2.49842453E+01                   4
C4H6O1-3OOH4            C   4H   7O   3    0G   300.000  5000.000 1386.000    41
 1.95456291E+01 1.60358540E-02-5.61768950E-06 8.86341914E-10-5.20072732E-14    2
-1.12679434E+04-6.99490153E+01 3.83045773E+00 5.07388403E-02-3.42226447E-05    3
 1.13486298E-08-1.48529245E-12-5.61786232E+03 1.51509867E+01                   4
C4H6O2-1OOH4            C   4H   7O   3    0G   300.000  5000.000 1364.000    41
 2.05164800E+01 1.55727845E-02-5.54197222E-06 8.83592649E-10-5.22241946E-14    2
-9.30030707E+03-7.46630628E+01 5.38344712E+00 4.47089832E-02-2.43630482E-05    3
 5.07835349E-09-1.20805939E-13-3.40711224E+03 8.84731441E+00                   4
HOCH2COCH2              C   3H   5O   2    0G   300.000  5000.000 1363.000    31
 1.27106963E+01 1.15513960E-02-3.95951917E-06 6.16237371E-10-3.58328248E-14    2
-2.71538154E+04-3.67129478E+01 4.98634970E+00 2.51766916E-02-1.10893306E-05    3
 1.12011467E-09 2.89491135E-13-2.40047973E+04 6.38258616E+00                   4
HOCH2CO    9/25/15      C   2H   3O   2    0G   300.000  5000.000 1487.000    21
 9.43496508E+00 7.68897340E-03-2.74959280E-06 4.39772312E-10-2.60488233E-14    2
-2.29700136E+04-2.04618579E+01 5.12916864E+00 9.07172819E-03 6.49228146E-06    3
-8.56591893E-09 2.31070825E-12-2.06151607E+04 5.73007596E+00                   4
HOCHCHO    9/25/15      C   2H   3O   2    0G   300.000  5000.000 1680.000    21
 9.99251726E+00 7.77560619E-03-2.94238616E-06 4.90136333E-10-2.98979778E-14    2
-2.20440827E+04-2.73957153E+01 5.42856274E-01 2.95295948E-02-2.08315490E-05    3
 6.72777461E-09-8.06116446E-13-1.89378452E+04 2.31681075E+01                   4
PC3H4OH-3  9/25/15      C   3H   5O   1    0G   300.000  5000.000 1378.000    11
 1.15297558E+01 1.14381097E-02-4.04415495E-06 6.41949269E-10-3.78242456E-14    2
-3.45486444E+03-3.65385497E+01 4.06368169E-01 3.70231405E-02-2.72202689E-05    3
 1.05783475E-08-1.73632514E-12 5.27160824E+02 2.34781848E+01                   4
PC3H4OH-1  9/25/15      C   3H   5O   1    0G   300.000  5000.000 1403.000    21
 1.09468986E+01 1.04014540E-02-3.44082448E-06 5.22105632E-10-2.98049266E-14    2
 4.11530600E+03-3.11161699E+01 2.07150195E+00 3.50016810E-02-3.01922013E-05    3
 1.38467853E-08-2.55380109E-12 6.81914209E+03 1.51916605E+01                   4
CH3COCHOH  9/25/15      C   3H   5O   2    0G   300.000  5000.000 1378.000    31
 1.23884831E+01 1.23099892E-02-4.32263800E-06 6.83043939E-10-4.01192794E-14    2
-2.97609476E+04-3.85682589E+01 2.11183979E+00 3.32521318E-02-1.96834015E-05    3
 5.40736760E-09-5.32450556E-13-2.58545486E+04 1.77643465E+01                   4
SC2H2OH    9/25/15      C   2H   3O   1    0G   300.000  5000.000 1410.000    11
 7.99235139E+00 5.83109353E-03-1.89242965E-06 2.83129118E-10-1.59933287E-14    2
 9.51237374E+03-1.62058375E+01 1.63791895E+00 2.64968839E-02-2.74821415E-05    3
 1.43110557E-08-2.85794966E-12 1.11467016E+04 1.58714777E+01                   4
PC4H8OH-1               C   4H   9O   1    0G   300.000  5000.000 1392.000    41
 1.47813217E+01 1.89692972E-02-6.38671427E-06 9.81341181E-10-5.65332084E-14    2
-1.88487062E+04-4.98892364E+01 7.72566991E-01 5.00429367E-02-3.20163534E-05    3
 1.02913291E-08-1.30709217E-12-1.38421800E+04 2.58928300E+01                   4
PC4H8OH-3               C   4H   9O   1    0G   300.000  5000.000 1398.000    41
 1.45944628E+01 1.92223378E-02-6.48868808E-06 9.98309067E-10-5.75488987E-14    2
-1.52392636E+04-4.85127747E+01 2.21685429E+00 4.71340178E-02-3.04254756E-05    3
 1.03165429E-08-1.45043599E-12-1.08208508E+04 1.83497891E+01                   4
C4H7O1-4   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1388.000    21
 1.33251126E+01 1.65057558E-02-5.65235890E-06 8.78319847E-10-5.09914580E-14    2
 1.91281414E+03-4.28181479E+01 2.44895430E+00 3.69423519E-02-1.77510852E-05    3
 2.64537530E-09 2.43666218E-13 6.16385921E+03 1.73174889E+01                   4
PC4H8OH-4               C   4H   9O   1    0G   300.000  5000.000 1401.000    41
 1.41519859E+01 1.96439700E-02-6.64537615E-06 1.02402720E-09-5.91001981E-14    2
-1.56141213E+04-4.50604102E+01-6.95634735E-02 5.20263179E-02-3.44849029E-05    3
 1.17704221E-08-1.63047436E-12-1.06053581E+04 3.15909567E+01                   4
SC4H8OH-2               C   4H   9O   1    0G   300.000  5000.000 1395.000    41
 1.45514712E+01 1.92722299E-02-6.50955109E-06 1.00200009E-09-5.77830714E-14    2
-2.09909632E+04-4.82454428E+01 1.96361387E+00 4.77673982E-02-3.11652479E-05    3
 1.07498897E-08-1.54834306E-12-1.65000330E+04 1.97286755E+01                   4
CH2COHCO   9/25/15      C   3H   3O   2    0G   300.000  5000.000 1411.000    11
 1.31285142E+01 6.17948608E-03-1.93387986E-06 2.81892606E-10-1.56244314E-14    2
-1.93507932E+04-4.22958094E+01 1.24341370E+00 4.71484739E-02-5.44200189E-05    3
 2.95970356E-08-6.01447282E-12-1.65555219E+04 1.68301276E+01                   4
C4H72-2O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1390.000    31
 1.63301022E+01 1.60698895E-02-5.50238293E-06 8.55098973E-10-4.96517196E-14    2
-4.70039715E+03-5.78736400E+01 2.49537080E+00 4.75680882E-02-3.26452548E-05    3
 1.14069694E-08-1.61494862E-12 1.76383849E+02 1.67027189E+01                   4
C4H71-1O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1390.000    31
 1.63738534E+01 1.62685376E-02-5.62192103E-06 8.78982520E-10-5.12510706E-14    2
-1.06318473E+03-5.69005716E+01 2.02223104E+00 4.85577506E-02-3.30293697E-05    3
 1.13406677E-08-1.57078109E-12 4.04143594E+03 2.06106646E+01                   4
C4H71-2O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1394.000    31
 1.63565639E+01 1.61768136E-02-5.56610316E-06 8.67700997E-10-5.04886444E-14    2
-3.40245466E+03-5.75260769E+01 1.42459973E+00 5.20547601E-02-3.89440869E-05    3
 1.51726193E-08-2.42611664E-12 1.68854104E+03 2.23230947E+01                   4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
 1.14795375E+01 1.45881429E-02-4.88359380E-06 7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01 1.13614529E+00 3.68850655E-02-2.24073579E-05    3
 6.62398992E-09-7.32206246E-13-1.09273174E+04 2.24919343E+01                   4
PC4H8OH-2O2             C   4H   9O   3    0G   300.000  5000.000 1407.000    51
 1.90513685E+01 2.00624257E-02-6.76970282E-06 1.04136985E-09-6.00271674E-14    2
-3.65966815E+04-6.71202048E+01 1.97780900E+00 6.25692373E-02-4.76730210E-05    3
 1.90561997E-08-3.10596799E-12-3.09625439E+04 2.35880251E+01                   4
SC4H8OH-1O2             C   4H   9O   3    0G   300.000  5000.000 1405.000    51
 1.88547090E+01 2.02217653E-02-6.82328766E-06 1.04961552E-09-6.05032676E-14    2
-3.65721162E+04-6.59105449E+01 1.47037864E+00 6.38295256E-02-4.92333916E-05    3
 1.99704964E-08-3.30499356E-12-3.08602292E+04 2.63462505E+01                   4
C4H71-3OOCH3            C   5H  10O   2    0G   300.000  5000.000 1387.000    51
 2.12299326E+01 2.07003584E-02-6.99464238E-06 1.07836941E-09-6.22999849E-14    2
-1.85005682E+04-8.53499854E+01-5.42404662E-01 7.51511469E-02-6.00684679E-05    3
 2.49701271E-08-4.22319878E-12-1.13061371E+04 3.02981962E+01                   4
C4H72-1OOCH3            C   5H  10O   2    0G   300.000  5000.000 1382.000    51
 1.92914755E+01 2.34475159E-02-8.16713690E-06 1.28338262E-09-7.50837828E-14    2
-1.72688938E+04-7.16509708E+01 2.44675386E+00 6.21430218E-02-4.39326296E-05    3
 1.72567499E-08-2.94950711E-12-1.11431755E+04 1.94028997E+01                   4
C4H6                    C   4H   6    0    0G   300.000  5000.000 1388.000    11
 1.01064561E+01 1.46248415E-02-5.01373934E-06 7.79510645E-10-4.52675769E-14    2
 9.96133753E+03-2.97310638E+01 1.01356056E+00 3.35722771E-02-1.96279376E-05    3
 5.74803850E-09-6.75029065E-13 1.33956759E+04 1.99957382E+01                   4
C4H612            A 8/83C   4H   6    0    0G   300.000  5000.000 1374.000    11
 1.14059885E+01 1.31489843E-02-4.43542071E-06 6.83028825E-10-3.94289265E-14    2
 1.42427294E+04-3.69674067E+01 9.45515689E-01 3.46162239E-02-1.98590697E-05    3
 5.02139421E-09-3.67977164E-13 1.81439079E+04 2.02191143E+01                   4
C4H6-2            A 8/83C   4H   6    0    0G   300.000  5000.000 1377.000    21
 9.60305554E+00 1.48972169E-02-5.16751230E-06 8.09757170E-10-4.72817668E-14    2
 1.24831314E+04-2.87129792E+01 1.97152408E+00 2.76790997E-02-1.13396645E-05    3
 1.02970745E-09 2.75290944E-13 1.57283766E+04 1.42147356E+01                   4
C4H5-I            H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1
 0.10229092E+02 0.94850138E-02-0.90406445E-07-0.12596100E-08 0.24781468E-12    2
 0.34642812E+05-0.28564529E+02-0.19932900E-01 0.38005672E-01-0.27559450E-04    3
 0.77835551E-08 0.40209383E-12 0.37496223E+05 0.24394241E+02                   4
C4H5-N            H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1
 0.98501978E+01 0.10779008E-01-0.13672125E-05-0.77200535E-09 0.18366314E-12    2
 0.38840301E+05-0.26001846E+02 0.16305321E+00 0.39830137E-01-0.34000128E-04    3
 0.15147233E-07-0.24665825E-11 0.41429766E+05 0.23536163E+02                   4
C4H5              H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1  ! lumped C4H5-N
 0.98501978E+01 0.10779008E-01-0.13672125E-05-0.77200535E-09 0.18366314E-12    2
 0.38840301E+05-0.26001846E+02 0.16305321E+00 0.39830137E-01-0.34000128E-04    3
 0.15147233E-07-0.24665825E-11 0.41429766E+05 0.23536163E+02                   4
C4H5-2            H6W/94C   4H   5    0    0G   300.000  5000.000 1385.000    11
 1.03230828E+01 1.17625574E-02-4.00004665E-06 6.18727929E-10-3.58083530E-14    2
 3.25861413E+04-2.88794317E+01 2.31011292E+00 2.83747046E-02-1.63836755E-05    3
 4.46251967E-09-4.30510879E-13 3.55842945E+04 1.49105965E+01                   4
C4H4              H6W/94C   4H   4    0    0G   300.000  3000.00  1000.00      1
 0.66507092E+01 0.16129434E-01-0.71938875E-05 0.14981787E-08-0.11864110E-12    2
 0.31195992E+05-0.97952118E+01-0.19152479E+01 0.52750878E-01-0.71655944E-04    3
 0.55072423E-07-0.17286228E-10 0.32978504E+05 0.31419983E+02                   4
C4H3-I            AB1/93C   4H   3    0    0G   300.000  3000.00  1000.00      1
 0.90978165E+01 0.92207119E-02-0.33878441E-05 0.49160498E-09-0.14529780E-13    2
 0.56600574E+05-0.19802597E+02 0.20830412E+01 0.40834274E-01-0.62159685E-04    3
 0.51679358E-07-0.17029184E-10 0.58005129E+05 0.13617462E+02                   4
C4H3-N            H6W/94C   4H   3    0    0G   300.000  3000.00  1000.00      1
 0.54328279E+01 0.16860981E-01-0.94313109E-05 0.25703895E-08-0.27456309E-12    2
 0.61600680E+05-0.15673981E+01-0.31684113E+00 0.46912100E-01-0.68093810E-04    3
 0.53179921E-07-0.16523005E-10 0.62476199E+05 0.24622559E+02                   4
C4H3              H6W/94C   4H   3    0    0G   300.000  3000.00  1000.00      1  ! lumped C4H3-N
 0.54328279E+01 0.16860981E-01-0.94313109E-05 0.25703895E-08-0.27456309E-12    2
 0.61600680E+05-0.15673981E+01-0.31684113E+00 0.46912100E-01-0.68093810E-04    3
 0.53179921E-07-0.16523005E-10 0.62476199E+05 0.24622559E+02                   4
C4H2              D11/99C   4H   2    0    0G   300.000  3000.000 1000.        1
 0.91576328E+01 0.55430518E-02-0.13591604E-05 0.18780075E-10 0.23189536E-13    2
 0.52588039E+05-0.23711460E+02 0.10543978E+01 0.41626960E-01-0.65871784E-04    3
 0.53257075E-07-0.16683162E-10 0.54185211E+05 0.14866591E+02                   4
C4H6O25           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
 8.60658242E+00 2.08310051E-02-8.42229481E-06 1.56717640E-09-1.09391202E-13    2
-1.76177415E+04-2.32464750E+01 2.67053463E+00 4.92586420E-03 8.86967406E-05    3
-1.26219194E-07 5.23991321E-11-1.46572472E+04 1.45722395E+01-1.30831522E+04    4
C2H3CHOCH2              C   4H   6O   1    0G   300.000  5000.000 1431.000    11
 1.26762790E+01 1.40819509E-02-4.63473868E-06 7.01090838E-10-3.99438277E-14    2
-4.08065264E+03-4.22515995E+01-3.59388437E+00 5.79063450E-02-4.97163294E-05    3
 2.15818682E-08-3.69199072E-12 8.58852628E+02 4.28475443E+01                   4
FURAN             T03/97C   4H   4O   1    0G   200.000  6000.0    1000.0      1
 9.38935003E+00 1.40291241E-02-5.07755110E-06 8.24137332E-10-4.95319963E-14    2
-8.68241814E+03-2.79162920E+01 8.47469463E-01 1.31773796E-02 5.99735901E-05    3
-9.71562904E-08 4.22733796E-11-5.36785445E+03 2.14945172E+01-4.17166616E+03    4
C4H6O23           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
 8.60658242E+00 2.08310051E-02-8.42229481E-06 1.56717640E-09-1.09391202E-13    2
-1.32392815E+04-2.32464750E+01 2.67053463E+00 4.92586420E-03 8.86967406E-05    3
-1.26219194E-07 5.23991321E-11-1.02787872E+04 1.45722395E+01-1.30831522E+04    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
 1.39299886E+01 1.13228814E-02-3.87393567E-06 6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01 4.51553480E-01 4.37530418E-02-3.37273602E-05    3
 1.31111496E-08-2.04732021E-12 2.14943141E+03 2.40835867E+01                   4
H2C4O             120189H   2C   4O   1     G  0300.00   4000.00  1000.00      1
 0.01026888E+03 0.04896164E-01-0.04885081E-05-0.02708566E-08 0.05107013E-12    2
 0.02346903E+06-0.02815985E+03 0.04810971E+02 0.01313999E+00 0.09865073E-05    3
-0.06120720E-07 0.01640003E-10 0.02545803E+06 0.02113424E+02                   4
NC3H7CHO   8/12/15      C   4H   8O   1    0G   300.000  5000.000 1679.000    31
 1.19789345E+01 2.04894148E-02-7.24831619E-06 1.15561709E-09-6.84119824E-14    2
-3.09272130E+04-3.63929716E+01 1.24208539E+00 4.21277518E-02-2.13832135E-05    3
 4.22614614E-09-1.03710908E-13-2.71049353E+04 2.21567167E+01                   4
NC3H7CO                 C   4H   7O   1    0G   300.000  5000.000 1496.000    31
 1.34870098E+01 1.58626861E-02-5.41698905E-06 8.40508889E-10-4.87570090E-14    2
-1.30725285E+04-4.38634081E+01 2.63537828E+00 3.40368642E-02-1.24118988E-05    3
-1.17886666E-09 1.16488136E-12-8.65919992E+03 1.68407569E+01                   4
C3H6CHO-1               C   4H   7O   1    0G   300.000  5000.000 1538.000    31
 1.33449137E+01 1.59347421E-02-5.43143577E-06 8.41706117E-10-4.87847084E-14    2
-6.91281947E+03-4.19662475E+01 2.21483383E+00 3.54113290E-02-1.44082892E-05    3
 5.27605922E-11 8.95003230E-13-2.46482792E+03 2.00076022E+01                   4
C3H6CHO-2               C   4H   7O   1    0G   300.000  5000.000 1439.000    31
 1.27128605E+01 1.68632757E-02-5.83779932E-06 9.14059755E-10-5.33575736E-14    2
-8.50165835E+03-3.84620358E+01 4.01372834E+00 2.33173718E-02 5.72463585E-06    3
-1.27182841E-08 3.69912722E-12-4.16766399E+03 1.30545921E+01                   4
C3H6CHO-3               C   4H   7O   1    0G   300.000  5000.000 1678.000    31
 1.21729663E+01 1.80056550E-02-6.43783092E-06 1.03362049E-09-6.14850407E-14    2
-1.08642352E+04-3.80322250E+01 5.29001237E-01 4.30707499E-02-2.49474118E-05    3
 6.40934608E-09-5.27769846E-13-6.87667117E+03 2.48856420E+01                   4
SC3H5CHO                C   4H   6O   1    0G   300.000  5000.000 1396.000    21
 1.33892118E+01 1.39115420E-02-4.75820958E-06 7.38736618E-10-4.28606559E-14    2
-1.97917448E+04-4.60146004E+01 1.09372823E+00 4.43315368E-02-3.41918451E-05    3
 1.39369607E-08-2.33791460E-12-1.56745978E+04 1.94458467E+01                   4
SC3H5CO                 C   4H   5O   1    0G   300.000  5000.000 1396.000    11
 1.29925654E+01 1.22140721E-02-4.19305277E-06 6.52697685E-10-3.79407376E-14    2
-2.74782380E+03-4.51092470E+01 7.76401404E-01 4.26828436E-02-3.37881191E-05    3
 1.39128174E-08-2.33331638E-12 1.29903132E+03 1.98102013E+01                   4
C2H5COCH3  8/12/15      C   4H   8O   1    0G   300.000  5000.000 1454.000    31
 1.28183044E+01 1.79874386E-02-5.94194784E-06 9.01636365E-10-5.14993729E-14    2
-3.51711964E+04-4.11609193E+01 2.57048052E+00 3.51446793E-02-1.23849584E-05    3
-1.21280927E-09 1.16163555E-12-3.10194049E+04 1.61395232E+01                   4
C2H5COCH2               C   4H   7O   1    0G   300.000  5000.000 1396.000    31
 1.35979480E+01 1.57187785E-02-5.35200820E-06 8.28428039E-10-4.79645862E-14    2
-1.30111973E+04-4.46215708E+01 1.96643032E+00 4.10271409E-02-2.56193885E-05    3
 7.86244495E-09-9.26825962E-13-8.80149212E+03 1.84803948E+01                   4
CH2CH2COCH3             C   4H   7O   1    0G   300.000  5000.000 1392.000    31
 1.17915603E+01 1.70296457E-02-5.75444256E-06 8.86035114E-10-5.11070778E-14    2
-9.70683178E+03-3.25532787E+01 2.36191763E+00 3.50400641E-02-1.70487065E-05    3
 3.09070210E-09 2.80364847E-14-6.02754073E+03 1.95184512E+01                   4
CH3CHCOCH3              C   4H   7O   1    0G   300.000  5000.000 1438.000    31
 1.19651378E+01 1.63142163E-02-5.39879520E-06 8.20454677E-10-4.69197541E-14    2
-1.51990676E+04-3.30142593E+01 3.31082456E+00 2.83712402E-02-5.64603859E-06    3
-4.62626296E-09 1.82954207E-12-1.14602301E+04 1.62217415E+01                   4
C2H3COCH3               C   4H   6O   1    0G   300.000  5000.000 1390.000    21
 1.19989844E+01 1.52616304E-02-5.26018882E-06 8.20774274E-10-4.77834528E-14    2
-2.12170620E+04-3.71383523E+01 6.55910700E-01 4.19405303E-02-3.00269693E-05    3
 1.16578089E-08-1.92100897E-12-1.72216627E+04 2.38412293E+01                   4
CH3CHOOCOCH3            C   4H   7O   3    0G   300.000  5000.000 1411.000    41
 1.68056216E+01 1.70791389E-02-5.69439450E-06 8.68878944E-10-4.98008338E-14    2
-3.06718613E+04-5.51178960E+01 4.30171569E+00 4.62273591E-02-3.12564494E-05    3
 1.08627824E-08-1.51478379E-12-2.63732146E+04 1.19724375E+01                   4
CH2CHOOHCOCH3           C   4H   7O   3    0G   300.000  5000.000 1413.000    51
 1.78031394E+01 1.60286227E-02-5.38152372E-06 8.25242310E-10-4.74718968E-14    2
-2.30767899E+04-5.87370258E+01 4.45962223E+00 4.67200276E-02-3.15878907E-05    3
 1.06245787E-08-1.38857032E-12-1.84720686E+04 1.29655977E+01                   4
C2H5CHCO                C   4H   6O   1    0G   300.000  5000.000 1550.000    21
-2.04040652E+02 2.93466880E-01-1.15884523E-04 1.95253673E-08-1.19030791E-12    2
 8.27380036E+04 1.21233386E+03-2.28307043E+01 1.70978191E-01-3.53394379E-04    3
 2.78221616E-07-6.77325074E-11-1.04125457E+04 1.31232921E+02                   4
IC4H6Q2-II 9/ 8/14      C   4H   8O   4    0G   300.000  5000.000 1386.000    61
 2.50360805E+01 1.60230197E-02-5.70704966E-06 9.10412038E-10-5.38294659E-14    2
-2.84196401E+04-9.67186452E+01 2.16408482E-01 8.25572149E-02-7.64540445E-05    3
 3.58211787E-08-6.67718658E-12-2.05694845E+04 3.36943223E+01                   4
C5H10-1                 C   5H  10    0    0G   300.000  5000.000 1390.000    31
 1.43624894E+01 2.26076154E-02-7.70500843E-06 1.19329968E-09-6.91126022E-14    2
-9.99915627E+03-5.12512094E+01-1.65023816E-01 5.30727359E-02-3.10861587E-05    3
 8.92413402E-09-9.81619602E-13-4.57363143E+03 2.80570113E+01                   4
C5H81-3    9/ 8/14      C   5H   8    0    0G   300.000  5000.000 1385.000    21
 1.29945372E+01 1.92678312E-02-6.58966712E-06 1.02295969E-09-5.93441369E-14    2
 4.59040047E+03-4.35689825E+01 1.54882436E+00 4.15042709E-02-2.14359890E-05    3
 4.71145517E-09-2.42142508E-13 9.05636062E+03 1.95665910E+01                   4
C5H9O1-3   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1379.000    31
 1.78860333E+01 2.04837367E-02-7.16613461E-06 1.12948597E-09-6.62221468E-14    2
-4.33139568E+03-6.72851315E+01 2.49666166E+00 5.20326105E-02-3.09828268E-05    3
 9.02567482E-09-1.04311127E-12 1.54758549E+03 1.70868328E+01                   4
BC5H10     9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1389.000    31
 1.40426423E+01 2.27915348E-02-7.74902598E-06 1.19814522E-09-6.93127003E-14    2
-1.32160483E+04-5.14469569E+01 6.04882839E-01 4.96635256E-02-2.66571142E-05    3
 6.47312078E-09-4.84017883E-13-8.06312207E+03 2.23818263E+01                   4
CC5H9-A                 C   5H   9    0    0G   300.000  5000.000 1393.000    31
 1.38635892E+01 2.06362872E-02-7.05717373E-06 1.09539676E-09-6.35381849E-14    2
 1.36104251E+04-4.72507189E+01-6.78909715E-01 5.37496002E-02-3.61116825E-05    3
 1.28563411E-08-1.92155723E-12 1.87974429E+04 3.12403382E+01                   4
CC5H9-B    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1392.000    21
 1.35249511E+01 2.14363755E-02-7.35304116E-06 1.14368637E-09-6.64363518E-14    2
 5.41381916E+03-5.00302394E+01-6.91501860E-01 5.09804846E-02-2.96448293E-05    3
 8.28273022E-09-8.57575066E-13 1.07478467E+04 2.76711552E+01                   4
AC5H9O-C                C   5H   9O   1    0G   300.000  5000.000 1382.000    31
 1.76789601E+01 2.05915073E-02-7.18764438E-06 1.13116483E-09-6.62505034E-14    2
-6.25146818E+03-6.62131721E+01 2.04951318E+00 5.36584877E-02-3.35086710E-05    3
 1.06174235E-08-1.39224338E-12-3.85112518E+02 1.91077262E+01                   4
CC5H9O-B   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1377.000    31
 1.86974377E+01 1.84542537E-02-6.18682537E-06 9.48850967E-10-5.46203980E-14    2
-7.15897769E+03-7.26540429E+01 2.75614808E+00 5.20514036E-02-3.10966938E-05    3
 8.25895065E-09-6.59917121E-13-1.35162741E+03 1.40990119E+01                   4
AC5H10                  C   5H  10    0    0G   300.000  5000.000 1392.000    31
 1.41931279E+01 2.26551019E-02-7.70008627E-06 1.19031326E-09-6.88489604E-14    2
-1.19491010E+04-5.10688681E+01-5.39429136E-01 5.44489715E-02-3.32707895E-05    3
 1.03047694E-08-1.28363329E-12-6.53967251E+03 2.90349986E+01                   4
AC5H9-A2                C   5H   9    0    0G   300.000  5000.000 1385.000    21
 1.50019889E+01 1.95965428E-02-6.60205927E-06 1.01535593E-09-5.85454957E-14    2
 5.90081014E+03-5.54528992E+01-9.54047710E-01 5.50153471E-02-3.58307910E-05    3
 1.16444141E-08-1.49086833E-12 1.15959514E+04 3.08476806E+01                   4
AC5H9-C                 C   5H   9    0    0G   300.000  5000.000 1392.000    21
 1.37918110E+01 2.09644966E-02-7.13793293E-06 1.10480881E-09-6.39628018E-14    2
 5.09555600E+03-5.01391436E+01-8.41372657E-01 5.27157283E-02-3.27334707E-05    3
 1.01974035E-08-1.26084730E-12 1.04321036E+04 2.93316754E+01                   4
AC5H9-D                 C   5H   9    0    0G   300.000  5000.000 1393.000    31
 1.35607521E+01 2.07514878E-02-7.06608626E-06 1.09362345E-09-6.33083050E-14    2
 1.31896844E+04-4.48718988E+01-1.67398152E-01 5.09876974E-02-3.22615638E-05    3
 1.05911843E-08-1.43705463E-12 1.81792947E+04 2.95710715E+01                   4
TC4H8CHO   9/ 7/95 THERMC   5H   9O   1    0G   300.000  5000.000 1397.00     41
 1.79663933E+01 1.94207117E-02-6.67409451E-06 1.03969221E-09-6.04702651E-14    2
-1.33368585E+04-6.79819424E+01-9.58078294E-01 6.42003258E-02-4.70776827E-05    3
 1.75737698E-08-2.64896151E-12-6.86582501E+03 3.33781112E+01                   4
O2C4H8CHO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1395.00     51
 2.12629904E+01 2.14072282E-02-7.38342949E-06 1.15281523E-09-6.71508438E-14    2
-3.16854524E+04-7.99828703E+01 1.91847699E+00 6.67245869E-02-4.80871046E-05    3
 1.78588690E-08-2.71163880E-12-2.49837984E+04 2.38577867E+01                   4
O2HC4H8CO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1394.00     61
 2.38219630E+01 1.91411448E-02-6.67919154E-06 1.05127303E-09-6.15876805E-14    2
-3.23093973E+04-9.42580755E+01 1.82607262E+00 6.93466111E-02-4.93125140E-05    3
 1.69848340E-08-2.26117657E-12-2.46578311E+04 2.41167544E+01                   4
C6H101-5   4/12/13 THERMC   6H  10    0    0G   300.000  5000.000 1413.000    21
 1.60456030E+01 2.34774145E-02-7.85797929E-06 1.20200542E-09-6.90100029E-14    2
 2.11899382E+03-5.88452460E+01-1.01375402E+00 6.38242808E-02-4.40653860E-05    3
 1.58295163E-08-2.30830701E-12 7.94033696E+03 3.25056094E+01                   4
C6H9-A    12/ 5/12 THERMC   6H   9    0    0G   300.000  5000.000 1400.000    21
 1.70842767E+01 2.08842788E-02-7.14529004E-06 1.10943563E-09-6.43676989E-14    2
 2.01040204E+04-6.39326012E+01-2.66715213E+00 7.26196475E-02-6.05323920E-05    3
 2.66000571E-08-4.74613408E-12 2.64415017E+04 4.02220332E+01                   4
IC4H7CHO                C   5H   8O   1    0G   300.000  5000.000 1391.000    31
 1.59171638E+01 1.93357284E-02-6.70857943E-06 1.05155191E-09-6.14175906E-14    2
-2.16140735E+04-5.67616631E+01-1.20982776E+00 5.92603375E-02-4.26960089E-05    3
 1.60356164E-08-2.49347521E-12-1.56205327E+04 3.53137305E+01                   4
L-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
 0.12715182E+02 0.13839662E-01-0.43765440E-05 0.31541636E-09 0.46619026E-13    2
 0.57031148E+05-0.39464600E+02 0.29590225E+00 0.58053318E-01-0.67766756E-04    3
 0.43376762E-07-0.11418864E-10 0.60001371E+05 0.22318970E+02                   4
C-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
 0.13849209E+02 0.78807920E-02 0.18243836E-05-0.21169166E-08 0.37459977E-12    2
 0.47446340E+05-0.50404953E+02-0.30991268E+01 0.54030564E-01-0.40839004E-04    3
 0.10738837E-07 0.98078490E-12 0.52205711E+05 0.37415207E+02                   4
C6H3              H6W/94C   6H   3    0    0G   300.000  3000.00  1000.00      1
 0.58188343E+01 0.27933408E-01-0.17825427E-04 0.53702536E-08-0.61707627E-12    2
 0.85188250E+05-0.92147827E+00 0.11790619E+01 0.55547360E-01-0.73076168E-04    3
 0.52076736E-07-0.15046964E-10 0.85647312E+05 0.19179199E+02                   4
!C6H2              P 1/93C   6H   2    0    0G   300.000  3000.00  1000.00      1 !ARAMCO
! 0.13226281E+02 0.73904302E-02-0.22715381E-05 0.25875217E-09-0.55356741E-14    2
! 0.80565258E+05-0.41201176E+02-0.15932624E+01 0.80530145E-01-0.14800649E-03    3
! 0.13300031E-06-0.45332313E-10 0.83273227E+05 0.27980873E+02                   4
C6H6              G 6/01C   6H   6    0    0G   200.000  6000.000 1000.000     1
 1.10809576E+01 2.07176746E-02-7.52145991E-06 1.22320984E-09-7.36091279E-14    2
 4.30641035E+03-4.00413310E+01 5.04818632E-01 1.85020642E-02 7.38345881E-05    3
-1.18135741E-07 5.07210429E-11 8.55247913E+03 2.16412893E+01 9.96811598E+03    4
FULVENE                0C   6H   6    0    0G   200.000  5000.000 1000.00    0 1 !Burcat kik
 1.14345282E+01 1.99371432E-02-7.13567060E-06 1.14951842E-09-6.87263886E-14    2
 2.04411455E+04-3.86799524E+01 5.09714763E-01 2.58195980E-02 5.06504954E-05    3
-9.32593825E-08 4.15963672E-11 2.44318827E+04 2.30638077E+01 2.60142888E+04    4
C6H5OOH    3/26/ 9 THERMC   6H   6O   2    0G   300.000  5000.000 1404.000    21
 1.92317474E+01 1.63154699E-02-5.53448904E-06 8.55059974E-10-4.94583790E-14    2
-1.01971012E+04-7.61674471E+01-4.03105975E+00 7.96101888E-02-7.21655013E-05    3
 3.27610696E-08-5.85584239E-12-3.10973017E+03 4.54324978E+01                   4
C6H5OH                  H   6C   6O   1    0G   300.000  5000.000 1417.000    01 !RDB: New Phenol Data from ATcT
 1.65836066E+01 1.68031411E-02-5.68590569E-06 8.76720329E-10-5.06327756E-14    2
-1.91953162E+04-6.64184870E+01-4.62896828E+00 7.24191655E-02-6.16064842E-05    3
 2.63313091E-08-4.44982390E-12-1.25672730E+04 4.51325260E+01                   4
C6H5O phenyox ra  T11/10C  6.H  5.O  1.   0.G   200.000  6000.000 1000.        1 !Burcat kik
 1.39194640E+01 1.82692821E-02-6.66348032E-06 1.08703146E-09-6.55586708E-14    2
 1.01826410E+03-5.03399303E+01-3.13089926E-01 3.91633523E-02 2.25817444E-05    3
-6.76854803E-08 3.28002121E-11 5.67534849E+03 2.71661147E+01 7.40392398E+03    4
C6H4OH     4/ 9/ 9 THERMC   6H   5O   1    0G   300.000  5000.000 1402.000    11
 1.73187560E+01 1.36366984E-02-4.68316332E-06 7.29071204E-10-4.23805358E-14    2
 1.14990276E+04-6.89986593E+01-5.99875435E+00 8.59063379E-02-9.12525636E-05    3
 4.72275890E-08-9.35576749E-12 1.78621926E+04 4.99931427E+01                   4
C5H6              T 1/90C   5H   6    0    0G   200.000  6000.000 1000.        1 !ARAMCO
 0.99757848E+01 0.18905543E-01-0.68411461E-05 0.11099340E-08-0.66680236E-13    2
 0.11081693E+05-0.32209454E+02 0.86108957E+00 0.14804031E-01 0.72108895E-04    3
-0.11338055E-06 0.48689972E-10 0.14801755E+05 0.21353453E+02 0.16152485E+05    4
!C5H6              T 1/90C   5H   6    0    0G   200.000  6000.000 1000.        1 !Burcat kik
! 9.88465785E+00 1.89943852E-02-6.87485480E-06 1.11556894E-09-6.70255571E-14    2
! 7.14353103E+03-3.17238367E+01 9.77484017E-01 1.39109570E-02 7.36279225E-05    3
!-1.14340239E-07 4.88766069E-11 1.08333853E+04 2.08861411E+01 1.21907364E+04    4
C5H6                    C   5H   6          G    200.00   3500.00 1000.00      1   ! 1705
 1.27914695e+00 3.77288105e-02-2.09426525e-05 5.50583680e-09-5.53554405e-13    2
 1.40655989e+04 1.47486951e+01-4.86268110e+00 6.22961227e-02-5.77936208e-05    3
 3.00731490e-08-6.69538246e-12 1.52939645e+04 4.43794652e+01                   4
C5H6-L     2/ 5/ 9 THERMC   5H   6    0    0G   300.000  5000.000 1372.000    21
 1.29600892E+01 1.48953758E-02-5.23622902E-06 8.27916389E-10-4.86464523E-14    2
 2.38180800E+04-4.25312093E+01 3.58448213E+00 3.24459626E-02-1.70150991E-05    3
 4.22715914E-09-4.18452556E-13 2.76514681E+04 9.60644208E+00                   4
C5H7       1/22/ 9 WKM  C   5H   7    0    0G   300.000  5000.000 1377.000    31
 1.36630213E+01 1.68061358E-02-5.98746539E-06 9.55341072E-10-5.64951981E-14    2
 1.27238941E+04-5.46331286E+01-6.75118368E+00 6.06461693E-02-4.01260152E-05    3
 1.22051562E-08-1.33459844E-12 2.01365277E+04 5.62694938E+01                   4
C5H5OH     5/ 2/91 THE.MC   5H   6O   1    0G   300.000  5000.000 1398.000    11
 1.53433477E+01 1.50754059E-02-5.13553582E-06 7.95807816E-10-4.61311517E-14    2
-1.19645453E+04-5.85204430E+01-4.26822012E+00 6.62446749E-02-5.68494038E-05    3
 2.46858526E-08-4.26820696E-12-5.75581338E+03 4.47962850E+01                   4
C5H5O      5/16/90 THERMC   5H   5O   1    0G   300.000  5000.000 1392.000    01
 1.48322894E+01 1.40483376E-02-4.92302051E-06 7.77041219E-10-4.56103939E-14    2
 1.45523665E+04-5.73228191E+01-2.83112840E+00 5.67277287E-02-4.44757303E-05    3
 1.74924447E-08-2.76004847E-12 2.04992154E+04 3.69634411E+01                   4
C5H3O            TAK0905C   5H   3O   1    0G   300.000  3500.000 1500.00      1
 1.19961781E+01 1.34287065E-02-5.90045309E-06 1.22553862E-09-9.86114716E-14    2
 2.89592010E+04-4.07548249E+01-3.03242604E+00 5.43937201E-02-4.95018348E-05    3
 2.25523751E-08-4.10727920E-12 3.35644081E+04 3.78374823E+01                   4
CVCCJCVC   3/1/95  Z&B  C   5H   7    0    0G   300.000  5000.000 1388.000    21
 1.40879309E+01 1.62398907E-02-5.64768950E-06 8.86857524E-10-5.18698993E-14    2
 1.76798698E+04-5.13735038E+01-2.94595603E+00 5.68783623E-02-4.31336497E-05    3
 1.68169537E-08-2.67926433E-12 2.35156925E+04 3.98188778E+01                   4
CVCCVCCJ           Z&B  C   5H   7    0    0G   300.000  5000.000 1386.000    21
 1.47302883E+01 1.59030900E-02-5.57729508E-06 8.80604825E-10-5.16963733E-14    2
 1.74050791E+04-5.42670706E+01-1.60087476E+00 5.38764703E-02-3.96302225E-05    3
 1.49599474E-08-2.31995284E-12 2.31199746E+04 3.35492960E+01                   4
CVCCJCVCOH 10/6/95 Z&B  C   5H   7O   1    0G   300.000  5000.000 1397.000    31
 1.67465815E+01 1.58357240E-02-5.44954706E-06 8.49881387E-10-4.94743246E-14    2
-4.30972870E+03-6.19378748E+01-2.91175436E+00 6.69362484E-02-5.71603047E-05    3
 2.48753749E-08-4.33243894E-12 1.96441523E+03 4.17454344E+01                   4
HOCVCCVO   1/26/ 9 WKM  C   3H   4O   2    0G   300.000  5000.000 1413.000    21
 1.66505478E+01 6.11745137E-03-2.09080785E-06 3.24985683E-10-1.88875073E-14    2
-3.82179939E+04-6.36794754E+01-2.01837189E+00 6.26539783E-02-6.73359280E-05    3
 3.39430425E-08-6.48917648E-12-3.31367523E+04 3.18162860E+01                   4
CVCCVCCOH  1/23/ 9 WKM  C   5H   8O   1    0G   300.000  5000.000 1396.000    31
 1.63079670E+01 1.79957763E-02-6.03115896E-06 9.23992259E-10-5.31254053E-14    2
-1.58204603E+04-5.84137244E+01-5.31488384E-01 6.06983915E-02-4.81499862E-05    3
 2.00308244E-08-3.38987282E-12-1.03301302E+04 3.07961436E+01                   4
OC5H7O     1/22/ 9 WKM  C   5H   7O   2    0G   300.000  5000.000 1375.000    31
 1.65416953E+01 1.86677673E-02-6.44836048E-06 1.00787611E-09-5.87521858E-14    2
-2.82017168E+04-5.47258181E+01 4.88394767E+00 4.03401300E-02-1.97774150E-05    3
 3.68903501E-09-3.40202384E-14-2.35295942E+04 9.97070337E+00                   4
OC4H6O     1/23/ 9 WKM  C   4H   6O   2    0G   300.000  5000.000 1382.000    31
 1.41894774E+01 1.53345510E-02-5.24594862E-06 8.14655154E-10-4.72759368E-14    2
-4.10001835E+04-4.43771751E+01 4.21628848E+00 3.57422725E-02-2.04226185E-05    3
 5.63821367E-09-5.88888993E-13-3.72055911E+04 1.02814620E+01                   4
OC4H5O     1/23/ 9 WKM  C   4H   5O   2    0G   300.000  5000.000 1388.000    21
 1.32138775E+01 1.37339051E-02-4.62639517E-06 7.10941370E-10-4.09538499E-14    2
-2.16535271E+04-3.64185255E+01 4.60550978E+00 3.30498712E-02-2.13102363E-05    3
 7.37021089E-09-1.08289438E-12-1.85460831E+04 1.01599453E+01                   4
O2CCHOOJ           Z&B  C   2H   1O   4    0G   300.000  5000.000 1682.000    01
 1.09910849E+01 7.46985861E-03-2.75568271E-06 4.51353051E-10-2.72108652E-14    2
-3.51335323E+04-2.11652231E+01 8.91497688E+00 8.60571847E-03 5.24416766E-07    3
-2.79301331E-09 7.62963051E-13-3.40867754E+04-8.72978273E+00                   4
HOCVCCJVO  1/26/ 9 WKM  C   3H   3O   2    0G   300.000  5000.000 1414.000    11
 1.52720985E+01 5.02586331E-03-1.68408578E-06 2.58390706E-10-1.48849424E-14    2
-1.98506828E+04-5.54641734E+01 6.07270082E-01 4.96011303E-02-5.32300885E-05    3
 2.68392951E-08-5.13094510E-12-1.58814562E+04 1.94817133E+01                   4
CJVCCVCCVO 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1396.000    21
 1.62360823E+01 1.18297101E-02-4.11454219E-06 6.46026823E-10-3.77767639E-14    2
 1.93499885E+04-5.83498817E+01-5.06628841E-01 6.04671965E-02-5.97396749E-05    3
 2.96804228E-08-5.76240010E-12 2.42765544E+04 2.82994148E+01                   4
CVCCVCCJVO 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1399.000    11
 1.53178248E+01 1.27352911E-02-4.35882964E-06 6.76912763E-10-3.92771371E-14    2
 7.60582726E+03-5.43599625E+01-2.18492198E-01 5.92100223E-02-5.89241174E-05    3
 2.97411920E-08-5.85244770E-12 1.20600764E+04 2.55968530E+01                   4
CJVCCVO    4/ 8/94 THERMC   3H   3O   1    0G   300.000  5000.000 1402.000    11
 1.07482537E+01 6.19822688E-03-2.06130981E-06 3.14418872E-10-1.80309517E-14    2
 1.51410162E+04-3.01266033E+01 1.46654466E+00 3.23390476E-02-3.05588208E-05    3
 1.44081861E-08-2.65600505E-12 1.78850058E+04 1.80850321E+01                   4
C#CCVCCJ           GLAR C   5H   5    0    0G   300.000  5000.000 1396.000    11
 1.41230912E+01 1.14233190E-02-3.95851276E-06 6.20128961E-10-3.62097887E-14    2
 4.25158384E+04-5.02942871E+01-6.16143558E-01 5.06466579E-02-4.48561743E-05    3
 2.02459419E-08-3.64542145E-12 4.71532377E+04 2.71623299E+01                   4
P-C6H3O2          AK0505C   6H   3O   2    0G   270.000  3000.000 1290.00      1
 1.22963699E+01 2.15055142E-02-1.07516136E-05 2.57528163E-09-2.41023652E-13    2
 1.15428998E+04-3.72584002E+01-1.57852347E+00 6.55376473E-02-6.50308721E-05    3
 3.32026554E-08-6.86665555E-12 1.51750093E+04 3.31518638E+01                   4
H15DE25DM               C   8H  14    0    0G   300.000  5000.000 1395.000    51
 2.25355644E+01 3.23955734E-02-1.10270814E-05 1.70640907E-09-9.87758061E-14    2
-1.04808866E+04-9.19784905E+01-1.71853441E+00 8.82613783E-02-6.03140500E-05    3
 2.15862289E-08-3.19690882E-12-1.95255748E+03 3.86048681E+01                   4
H15DE25DM-S             C   8H  13    0    0G   300.000  5000.000 1395.000    41
 2.21422958E+01 3.06966055E-02-1.04617380E-05 1.62037747E-09-9.38578511E-14    2
 6.56045671E+03-9.04059585E+01-2.04235551E+00 8.66261688E-02-5.99110976E-05    3
 2.15551630E-08-3.18976697E-12 1.50224279E+04 3.96917763E+01                   4
H15DE25DM-A             C   8H  13    0    0G   300.000  5000.000 1391.000    41
 2.33282646E+01 2.93694154E-02-9.94258906E-06 1.53368063E-09-8.86030202E-14    2
 7.37319036E+03-9.55902415E+01-2.21863377E+00 8.91652629E-02-6.33360636E-05    3
 2.32007379E-08-3.46329567E-12 1.61971179E+04 4.15116620E+01                   4
H15DE25DM-AO            C   8H  13O   1    0G   300.000  5000.000 1378.000    51
 2.50985951E+01 3.15085628E-02-1.10076915E-05 1.73332426E-09-1.01557468E-13    2
-2.49465338E+03-1.01097942E+02 3.03691957E+00 7.50640438E-02-4.17779534E-05    3
 1.07915725E-08-9.97734397E-13 6.11649780E+03 2.04746031E+01                   4
H15DE25DM-SO            C   8H  13O   1    0G   300.000  5000.000 1388.000    51
 2.60152179E+01 3.04295766E-02-1.05676513E-05 1.65746547E-09-9.68470091E-14    2
-4.79568520E+03-1.06442472E+02 9.30464015E-01 8.71669873E-02-5.99582593E-05    3
 2.15026041E-08-3.21687573E-12 4.19310073E+03 2.90924508E+01                   4
H15DE2M-T               C   7H  11    0    0G   300.000  5000.000 1389.000    41
 1.90144729E+01 2.61932198E-02-9.01183878E-06 1.40455988E-09-8.17075251E-14    2
 2.35551101E+04-7.15568628E+01 3.88856066E-01 6.70215700E-02-4.29671268E-05    3
 1.42489875E-08-1.96105571E-12 3.03627273E+04 2.95444186E+01                   4
B2E2M1OJ                C   5H   9O   1    0G   300.000  5000.000 2003.000    31
 1.35666458E+01 2.56547934E-02-9.37226256E-06 1.52518398E-09-9.15378763E-14    2
-3.58767067E+03-4.27272791E+01 5.64762692E+00 3.43609862E-02-5.60649548E-06    3
-5.19111402E-09 1.73155461E-12-6.65737793E+00 3.13825267E+00                   4
B13DE2M                 C   5H   8    0    0G   300.000  5000.000 1397.000    21
 1.40757545E+01 1.82375566E-02-6.20747687E-06 9.60350919E-10-5.55741525E-14    2
 2.40033881E+03-5.12988284E+01-4.72170009E-01 5.59413257E-02-4.50458826E-05    3
 1.96181377E-08-3.52009647E-12 7.14960489E+03 2.56276807E+01                   4
B13DE2MJ                C   5H   7    0    0G   300.000  5000.000 1393.000    11
 1.48413344E+01 1.52425753E-02-5.13559858E-06 7.89787260E-10-4.55353492E-14    2
 2.02661570E+04-5.54474955E+01-8.98037227E-01 5.65174321E-02-4.76107829E-05    3
 2.09672106E-08-3.73076319E-12 2.52881763E+04 2.74966602E+01                   4
B12DE3M   11/12/12 THERMC   5H   8    0    0G   300.000  5000.000 1388.000    21
 1.37093177E+01 1.85726726E-02-6.33115904E-06 9.80719059E-10-5.68099894E-14    2
 8.59518752E+03-4.88749621E+01 1.27860173E+00 4.54917474E-02-2.82334169E-05    3
 8.98449372E-09-1.17220042E-12 1.31637341E+04 1.87039373E+01                   4
B2E3M1OJ                C   5H   9O   1    0G   300.000  5000.000 2003.000    31
 1.35666458E+01 2.56547934E-02-9.37226256E-06 1.52518398E-09-9.15378763E-14    2
-3.58767067E+03-4.27272791E+01 5.64762692E+00 3.43609862E-02-5.60649548E-06    3
-5.19111402E-09 1.73155461E-12-6.65737793E+00 3.13825267E+00                   4
C8H141-5,3-4            C   8H  14    0    0G   300.000  5000.000 1396.000    51
 2.30690680E+01 3.23154042E-02-1.10795683E-05 1.72276354E-09-1.00052582E-13    2
-8.91240214E+03-9.49655754E+01-2.52713194E+00 9.28837673E-02-6.67176819E-05    3
 2.53683579E-08-4.01212661E-12-4.55965940E+01 4.23180878E+01                   4
C8H141-5,3  8/25/15     C   8H  14    0    0G   300.000  5000.000 1392.000    51
 2.25173982E+01 3.26748629E-02-1.11807923E-05 1.73629966E-09-1.00752481E-13    2
-8.96062790E+03-9.10857551E+01-1.02072126E+00 8.47808555E-02-5.47568199E-05    3
 1.81792070E-08-2.47335881E-12-4.53248586E+02 3.64247438E+01                   4
C8H142-6   8/25/15      C   8H  14    0    0G   300.000  5000.000 1386.000    51
 2.20960852E+01 3.27887472E-02-1.11700037E-05 1.72970378E-09-1.00179059E-13    2
-9.04951881E+03-8.92942652E+01 3.43524821E-01 7.72359120E-02-4.34861460E-05    3
 1.12949093E-08-9.77995416E-13-8.37798357E+02 2.98241439E+01                   4
C8H131-5,3-4,TA         C   8H  13    0    0G   300.000  5000.000 1394.000    41
 2.22822575E+01 3.10651867E-02-1.06940907E-05 1.66739777E-09-9.70243450E-14    2
 7.57680613E+03-9.19858764E+01-3.23996819E+00 9.13494930E-02-6.60037456E-05    3
 2.51706078E-08-3.99030974E-12 1.64345368E+04 4.49498860E+01                   4
C8H131-5,3,TA           C   8H  13    0    0G   300.000  5000.000 1389.000    41
 2.16161787E+01 3.14326704E-02-1.07786324E-05 1.67632587E-09-9.73755313E-14    2
 7.60897211E+03-8.80384104E+01-5.03201172E-01 7.78854227E-02-4.63156182E-05    3
 1.32834166E-08-1.42623050E-12 1.58388712E+04 3.26514434E+01                   4
C8H131-5,3,SA           C   8H  13    0    0G   300.000  5000.000 1392.000    41
 2.21141889E+01 3.09871348E-02-1.06198459E-05 1.65100088E-09-9.58788408E-14    2
 8.08509780E+03-9.01448021E+01-1.32185914E+00 8.30473789E-02-5.42213233E-05    3
 1.80737386E-08-2.45105483E-12 1.65183103E+04 3.67169651E+01                   4
C8H131-5,3,PA           C   8H  13    0    0G   300.000  5000.000 1389.000    41
 2.32085707E+01 2.97529224E-02-1.01333635E-05 1.56925634E-09-9.09001242E-14    2
 8.95338901E+03-9.40777602E+01-1.57063382E+00 8.60080913E-02-5.83884368E-05    3
 2.02048105E-08-2.83115953E-12 1.77015232E+04 3.95476224E+01                   4
C8H132-6,SA             C   8H  13    0    0G   300.000  5000.000 1387.000    41
 2.16167233E+01 3.12260643E-02-1.06640216E-05 1.65409816E-09-9.59112187E-14    2
 8.03384556E+03-8.72194430E+01 2.20017932E-01 7.48621425E-02-4.21239973E-05    3
 1.07414215E-08-8.66560315E-13 1.61027987E+04 2.99517204E+01                   4
C8H132-6,PA             C   8H  13    0    0G   300.000  5000.000 1378.000    41
 2.29293875E+01 2.97187394E-02-1.00712335E-05 1.55505094E-09-8.99129602E-14    2
 8.77975921E+03-9.24517461E+01 1.05119796E-01 7.70150350E-02-4.48890925E-05    3
 1.19516688E-08-1.04377517E-12 1.72713386E+04 3.22058738E+01                   4
C6H101-3,3              C   6H  10    0    0G   300.000  5000.000 1395.000    31
 1.69678361E+01 2.28868236E-02-7.78758381E-06 1.20465198E-09-6.97080856E-14    2
-2.97276905E+03-6.58632941E+01-3.01310455E-02 6.43105079E-02-4.75083462E-05    3
 1.89877768E-08-3.17681035E-12 2.82367411E+03 2.49254708E+01                   4
C8H131-5,3-4,TAO        C   8H  13O   1    0G   300.000  5000.000 1394.000    51
 2.70579050E+01 2.84726632E-02-9.66434779E-06 1.49337149E-09-8.63788413E-14    2
-4.43111126E+03-1.12228392E+02 1.00679908E+00 8.90191278E-02-6.27963646E-05    3
 2.24161585E-08-3.20587060E-12 4.56422741E+03 2.76546640E+01                   4
C8H131-5,3,TAO          C   8H  13O   1    0G   300.000  5000.000 1396.000    51
 2.16638860E+01 2.77253448E-02-9.69375951E-06 1.67582120E-09-1.08059396E-13    2
-5.70300683E+03-9.33237797E+01 1.46771925E+00 7.67800622E-02-5.63189881E-05    3
 2.22689786E-08-3.64813515E-12 1.17475936E+03 1.45619856E+01                   4
C8H131-5,3,SAO          C   8H  13O   1    0G   300.000  5000.000 1385.000    51
 2.61023602E+01 3.05036647E-02-1.06268215E-05 1.67026867E-09-9.77389024E-14    2
-3.64744193E+03-1.06781316E+02 1.60953926E+00 8.39738786E-02-5.49469234E-05    3
 1.84255257E-08-2.56040058E-12 5.33713436E+03 2.62653941E+01                   4
C8H131-5,3,PAO          C   8H  13O   1    0G   300.000  5000.000 1374.000    51
 2.51902631E+01 3.15630048E-02-1.10568300E-05 1.74424175E-09-1.02327221E-13    2
-1.34401684E+03-1.01448477E+02 3.91532442E+00 7.10319966E-02-3.55623644E-05    3
 6.98595095E-09-1.83465840E-13 7.22911524E+03 1.67145758E+01                   4
C8H132-6,SAO            C   8H  13O   1    0G   300.000  5000.000 1381.000    51
 2.54267504E+01 3.10421548E-02-1.08045689E-05 1.69716523E-09-9.92701997E-14    2
-3.28641768E+03-1.02872762E+02 3.34168622E+00 7.49917518E-02-4.18382842E-05    3
 1.06108028E-08-8.96488454E-13 5.24458399E+03 1.86128166E+01                   4
C8H132-6,PAO            C   8H  13O   1    0G   300.000  5000.000 2014.000    51
 1.99391776E+01 3.79081645E-02-1.37893231E-05 2.23770591E-09-1.34044177E-13    2
 1.42981257E+03-7.07923233E+01 6.30807632E+00 5.80374259E-02-1.75637726E-05    3
-2.70887760E-09 1.61702129E-12 7.07839485E+03 6.29344560E+00                   4
C7H111-5,3,6P           C   7H  11    0    0G   300.000  5000.000 1396.000    41
 1.95787047E+01 2.54213538E-02-8.68127275E-06 1.34629701E-09-7.80464853E-14    2
 2.58537943E+04-7.44112330E+01-6.76848821E-01 7.38082653E-02-5.35945220E-05    3
 2.06293915E-08-3.29701110E-12 3.28160434E+04 3.40518079E+01                   4
C7H111-5,1P             C   7H  11    0    0G   300.000  5000.000 1388.000    41
 1.91915682E+01 2.55013021E-02-8.65881522E-06 1.33796943E-09-7.73784878E-14    2
 2.60946287E+04-7.21387547E+01 8.16831855E-01 6.56745024E-02-4.14490949E-05    3
 1.32234876E-08-1.69289568E-12 3.27646149E+04 2.75442934E+01                   4
C4H64,2-1OH             C   4H   7O   1    0G   300.000  5000.000 1366.000    21
 1.36259446E+01 1.70233137E-02-6.00460246E-06 9.51603754E-10-5.60055773E-14    2
-7.81498890E+03-4.44948073E+01 2.50804582E+00 3.53393033E-02-1.41418095E-05    3
 5.65501810E-10 5.94838384E-13-3.08574102E+03 1.81061546E+01                   4
C4H63,1-1OH             C   4H   7O   1    0G   300.000  5000.000 1401.000    21
 1.38675222E+01 1.54795810E-02-5.17720236E-06 7.91828077E-10-4.54656891E-14    2
-1.07655481E+04-4.87820652E+01-5.96640682E-01 5.31885124E-02-4.34791765E-05    3
 1.86514084E-08-3.23780972E-12-6.15543596E+03 2.74734171E+01                   4
C4H63,1-3OH             C   4H   7O   1    0G   300.000  5000.000 1380.000    21
 1.33633351E+01 1.70222596E-02-5.95245190E-06 9.37896168E-10-5.49767305E-14    2
-9.90113178E+03-4.54753472E+01 5.96155469E-01 4.35893351E-02-2.65985265E-05    3
 8.14250262E-09-1.02316366E-12-5.05630797E+03 2.43923636E+01                   4
C4H63,1-2OH             C   4H   7O   1    0G   300.000  5000.000 1404.000    21
 1.46899596E+01 1.48008021E-02-4.94483770E-06 7.55542892E-10-4.33461574E-14    2
-1.29448240E+04-5.45653093E+01-1.58903600E+00 6.17722944E-02-5.78263835E-05    3
 2.78090017E-08-5.26779799E-12-8.17977186E+03 2.96999338E+01                   4
C4H5OH-13  9/24/15      C   4H   6O   1    0G   300.000  5000.000 1405.000    21
 1.40975061E+01 1.29826578E-02-4.36356696E-06 6.69260196E-10-3.84920001E-14    2
-1.41099189E+04-4.94340793E+01-1.60022758E+00 6.12386329E-02-6.18933585E-05    3
 3.14927455E-08-6.20396658E-12-9.77435172E+03 3.08328186E+01                   4
SQC4H7OHP-4             C   4H   9O   3    0G   300.000  5000.000 1410.000    61
 1.99207495E+01 1.89422879E-02-6.39488327E-06 9.84231371E-10-5.67606301E-14    2
-2.89250584E+04-7.01061222E+01 1.44518283E+00 6.52944119E-02-5.10380130E-05    3
 2.05238910E-08-3.32050656E-12-2.29059890E+04 2.78546218E+01                   4
CY(CCCO)COH             C   4H   8O   2    0G   300.000  5000.000 1396.000    21
 1.34636332E+01 2.28745777E-02-9.93619553E-06 1.89605197E-09-1.26466856E-13    2
-3.96396606E+04-4.51064489E+01-6.97589766E+00 7.98392838E-02-7.11131714E-05    3
 3.16611877E-08-5.61324136E-12-3.35777839E+04 6.12093340E+01                   4
SQC4H7OHP-4O2           C   4H   9O   5    0G   300.000  5000.000 1402.000    71
 2.35936348E+01 2.08588461E-02-7.13602285E-06 1.10820581E-09-6.43133049E-14    2
-4.78452356E+04-8.49505816E+01 2.62618431E+00 7.26812595E-02-5.64956508E-05    3
 2.25892409E-08-3.65246549E-12-4.08999596E+04 2.65615323E+01                   4
PQC4H7OHS-3O2           C   4H   9O   5    0G   300.000  5000.000 1414.000    71
 2.46607662E+01 1.92947770E-02-6.45433722E-06 9.87246207E-10-5.66889630E-14    2
-4.98467067E+04-9.10424907E+01 2.90986916E+00 7.76596028E-02-6.68513896E-05    3
 2.93627835E-08-5.12008013E-12-4.31551961E+04 2.29130715E+01                   4
SQC4H7OHS-4O2           C   4H   9O   5    0G   300.000  5000.000 1414.000    71
 2.46607662E+01 1.92947770E-02-6.45433722E-06 9.87246207E-10-5.66889630E-14    2
-4.98467067E+04-9.10424907E+01 2.90986916E+00 7.76596028E-02-6.68513896E-05    3
 2.93627835E-08-5.12008013E-12-4.31551961E+04 2.29130715E+01                   4
C4H7O2-1,3OOH           C   4H   9O   5    0G   300.000  5000.000 1425.000    71
 2.54691227E+01 1.86441036E-02-6.23825706E-06 9.54422873E-10-5.48154425E-14    2
-4.01531561E+04-9.60389710E+01 4.88339443E+00 7.18219147E-02-5.86792171E-05    3
 2.42823866E-08-3.98538527E-12-3.36575518E+04 1.24696185E+01                   4
SC4H8OH-3O2             C   4H   9O   3    0G   300.000  5000.000 1417.000    51
 1.93082953E+01 1.92156764E-02-6.34250732E-06 9.60912935E-10-5.47939937E-14    2
-3.84370805E+04-6.88887622E+01 1.78918281E+00 6.62988026E-02-5.52280656E-05    3
 2.40247962E-08-4.18762027E-12-3.30428157E+04 2.28885942E+01                   4
CCY(COCC)OH             C   4H   8O   2    0G   300.000  5000.000 1328.000    21
 1.03816782E+01 2.53052690E-02-1.00511826E-05 1.68204740E-09-9.58092966E-14    2
-3.94348914E+04-2.73522595E+01-6.13260697E+00 7.75376285E-02-6.73066149E-05    3
 2.82841623E-08-4.65470382E-12-3.57825027E+04 5.53089299E+01                   4
COHQCYC(COC)            C   4H   8O   4    0G   300.000  5000.000 1319.000    51
 2.44599226E+01 1.64187782E-02-5.74024372E-06 9.05710407E-10-5.31829152E-14    2
-6.01811228E+04-1.02049722E+02 2.40687943E+00 5.95180442E-02-3.16913659E-05    3
 4.23694824E-09 8.42033474E-13-5.19694864E+04 1.88941416E+01                   4
QCYC(CCOC)OH            C   4H   8O   4    0G   300.000  5000.000 1411.000    41
 2.20860197E+01 1.83743733E-02-6.29478769E-06 9.78787994E-10-5.68621317E-14    2
-5.89652037E+04-8.64964494E+01-2.09099972E+00 8.02656739E-02-6.69756245E-05    3
 2.79282034E-08-4.60981823E-12-5.12529252E+04 4.11897260E+01                   4
HOCOCQ(CH3)2            C   4H   8O   4    0G   300.000  5000.000 1380.000    61
 2.28935401E+01 1.78627606E-02-6.34627520E-06 1.01068546E-09-5.96885712E-14    2
-8.05400680E+04-9.08953779E+01 1.56326363E+00 6.77165643E-02-5.14600149E-05    3
 1.99184629E-08-3.16007445E-12-7.30943302E+04 2.37255421E+01                   4
IQC4H7OHTO2             C   4H   9O   5    0G   300.000  5000.000 1389.000    71
 2.41720261E+01 2.09397176E-02-7.29061406E-06 1.14554056E-09-6.70217517E-14    2
-5.04772118E+04-8.95996685E+01 3.83287364E+00 6.90926177E-02-5.15031144E-05    3
 1.99235553E-08-3.17456897E-12-4.34442789E+04 1.94648622E+01                   4
IQC4H8OTQ-I             C   4H   9O   5    0G   300.000  5000.000 1386.000    71
 2.53249383E+01 2.00634820E-02-7.01249558E-06 1.10475030E-09-6.47561724E-14    2
-4.09610593E+04-9.73592779E+01 5.90219800E+00 6.26952142E-02-4.17351838E-05    3
 1.35422162E-08-1.71169663E-12-3.39620020E+04 7.89290087E+00                   4
IQC4H7OHTQ-P            C   4H   9O   5    0G   300.000  5000.000 1391.000    81
 2.45769593E+01 2.01889393E-02-7.03584537E-06 1.10623327E-09-6.47523225E-14    2
-4.25783112E+04-9.05052742E+01 3.45242802E+00 7.14541224E-02-5.54616790E-05    3
 2.22754676E-08-3.66067450E-12-3.54133076E+04 2.23024492E+01                   4
CHOC(CH3)OHCH2Q         C   4H   8O   4    0G   300.000  5000.000 1383.000    61
 2.24480753E+01 1.78753902E-02-6.26904597E-06 9.90084046E-10-5.81417382E-14    2
-6.55093075E+04-8.56747327E+01 2.40933530E+00 6.13326038E-02-4.03874986E-05    3
 1.22738404E-08-1.32997480E-12-5.83049516E+04 2.29870742E+01                   4
CO(CH2OOH)2             C   3H   6O   5    0G   300.000  5000.000 1393.000    61
 2.43376341E+01 1.14074110E-02-4.08931881E-06 6.55183244E-10-3.88570518E-14    2
-5.16862647E+04-9.01518175E+01-2.47626577E+00 8.93736793E-02-9.25891121E-05    3
 4.63168490E-08-8.93300309E-12-4.38924057E+04 4.84479477E+01                   4
AR                G 5/97AR  1  0    0      0G   200.000  6000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 4.37967491E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 4.37967491E+00 0.00000000E+00    4
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2
-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3
 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00 0.00000000E+00    4
HE                G 5/97HE 1    0    0    0 G   200.000  6000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 9.28723974E-01 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 9.28723974E-01 0.00000000E+00    4
IC3H7      8/12/15      C   3H   7    0    0G   298.000  5000.000 1000.000    21  
 6.70775549E+00 1.74048076E-02-6.07615926E-06 9.60084351E-10-5.65656490E-14    2
 7.55377821E+03-1.03686516E+01-8.97467137E-01 4.15744022E-02-4.94778349E-05    3
 4.56493655E-08-1.79085437E-11 9.93950407E+03 2.92641758E+01                   4
NC3H7      8/12/15      C   3H   7    0    0G   298.000  5000.000 1000.000    21
 7.48614243E+00 1.65769478E-02-5.74876481E-06 9.04103694E-10-5.30867231E-14    2
 8.93710008E+03-1.42595379E+01-2.20120865E+00 5.29641653E-02-7.23640506E-05    3
 6.36996940E-08-2.29332581E-11 1.15130744E+04 3.43669174E+01                   4
BIN1A                   C  20H  16          G   300.00   4000.00  1000.00      1
 .384004130e+02 .613760802e-01-.226838420e-04 .377828116e-08-.235041851e-12    2
-.165747108e+04-.190858878e+03-.946290891e+01 .179252381e+00-.989756752e-04    3
-.116559979e-07 .214782048e-10 .122142317e+05 .597553003e+02                   4
BIN1B                   C  20H  10          G   300.00   4000.00  1000.00      1
 .329670254e+02 .526917977e-01-.194742383e-04 .324368101e-08-.201785086e-12    2
 .107718330e+04-.161481167e+03-.895697031e+01 .146820540e+00-.577692501e-04    3
-.392441219e-07 .283752285e-10 .136083600e+05 .601566475e+02                   4
BIN1C                   C  20H   5          G   300.00   4000.00  1000.00      1
 .288518394e+02 .461144212e-01-.170433212e-04 .283878100e-08-.176596796e-12    2
-.612310898e+04-.152441597e+03-.829114243e+01 .126981825e+00-.389276128e-04    3
-.485387475e-07 .293596977e-10 .481805809e+04 .439495435e+02                   4
BIN2A                   C  40H  31          G   300.00   4000.00  1000.00      1
 .759883346e+02 .121453540e+00-.448877300e-04 .747661988e-08-.465110589e-12    2
 .397395323e+03-.376351286e+03-.224069955e+02 .373191638e+00-.228373343e-03    3
 .179614865e-08 .353583380e-10 .283409758e+05 .136281912e+03                   4
BIN2B                   C  40H  16          G   300.00   4000.00  1000.00      1
 .626025956e+02 .100058870e+00-.369805239e-04 .615957460e-08-.383178953e-12    2
-.435148944e+04-.314195266e+03-.175541017e+02 .277427018e+00-.990102332e-04    3
-.875044514e-07 .580969283e-10 .195176885e+05 .109755604e+03                   4
BIN2C                   C  40H   8          G   300.00   4000.00  1000.00      1
 .559396852e+02 .894094194e-01-.330446185e-04 .550399973e-08-.342396515e-12    2
-.170085815e+05-.296661132e+03-.168344238e+02 .244998896e+00-.659536990e-04    3
-.105536867e-06 .607898710e-10 .447424565e+04 .886402226e+02                   4
BIN3A                   C  80H  60          G   300.00   4000.00  1000.00      1
 .150797478e+03 .241022357e+00-.890788896e-04 .148372172e-07-.923003567e-12    2
 .303189596e+04-.764406699e+03-.455633619e+02 .756332498e+00-.489114578e-03    3
 .351844886e-07 .598168799e-10 .578481001e+05 .254746237e+03                   4
BIN3B                   C  80H  24          G   300.00   4000.00  1000.00      1
 .118542281e+03 .189468289e+00-.700251424e-04 .116635743e-07-.725575467e-12    2
-.213600710e+05-.610856398e+03-.343885254e+02 .522425915e+00-.164963932e-03    3
-.193041318e-06 .118886799e-09 .239919342e+05 .198395827e+03                   4
BIN3C                   C  80H   8          G   300.00   4000.00  1000.00      1
 .105216460e+03 .168169388e+00-.621533316e-04 .103524246e-07-.644010591e-12    2
-.466742552e+05-.575788129e+03-.329491696e+02 .457569671e+00-.988508639e-04    3
-.229106149e-06 .124272685e-09-.609495158e+04 .156165064e+03                   4
BIN4A                   C 160H 116          G   300.00   4000.00  1000.00      1
 .299236573e+03 .478275269e+00-.176764639e-03 .294423892e-07-.183157191e-11    2
 .105380025e+05-.155222165e+04-.926254655e+02 .153256344e+01-.104296494e-02    3
 .133553360e-06 .978341677e-10 .118028497e+06 .473857298e+03                   4
BIN4B                   C 160H  32          G   300.00   4000.00  1000.00      1
 .223758741e+03 .357637678e+00-.132178474e-03 .220159989e-07-.136958606e-11    2
-.680343262e+05-.118664453e+04-.673376950e+02 .979995585e+00-.263814796e-03    3
-.422147467e-06 .243159484e-09 .178969826e+05 .354560890e+03                   4
BIN4C                   C 160H  10          G   300.00   4000.00  1000.00      1
 .205435737e+03 .328351689e+00-.121354734e-03 .202131681e-07-.125743435e-11    2
-.102752674e+06-.113842566e+04-.653585808e+02 .890818250e+00-.172909327e-03    3
-.471736610e-06 .250565077e-09-.233838303e+05 .296493591e+03                   4
BIN5A                   C 320H 224          G   300.00   4000.00  1000.00      1
 .593310588e+03 .948299129e+00-.350479658e-03 .583768256e-07-.363154476e-11    2
 .352119959e+05-.312882274e+04-.194461399e+03 .312434830e+01-.224387754e-02    3
 .412099583e-06 .147772804e-09 .247380465e+06 .927804457e+03                   4
BIN5B                   C 320H  64          G   300.00   4000.00  1000.00      1
 .447517482e+03 .715275356e+00-.264356948e-03 .440319979e-07-.273917212e-11    2
-.135714032e+06-.237328905e+04-.134675390e+03 .195999117e+01-.527629592e-03    3
-.844294935e-06 .486318968e-09 .361485852e+05 .709121781e+03                   4
BIN5C                   C 320H  18          G   300.00   4000.00  1000.00      1
 .409205747e+03 .654041015e+00-.241725492e-03 .402624424e-07-.250467310e-11    2
-.208758277e+06-.227246778e+04-.130537242e+03 .177352947e+01-.337554521e-03    3
-.947981323e-06 .501803389e-09-.506171764e+05 .587708337e+03                   4
BIN6A                   C 640H 432          G   300.00   4000.00  1000.00      1
 .117696475e+04 .188116422e+01-.695255086e-03 .115803539e-06-.720398434e-11    2
 .909146192e+05-.634005997e+04-.398024258e+03 .633800264e+01-.476093625e-02    3
 .108624875e-05 .206199066e-09 .507419557e+06 .173874832e+04                   4
BIN6B                   C 640H 128          G   300.00   4000.00  1000.00      1
 .895034964e+03 .143055071e+01-.528713896e-03 .880639958e-07-.547834423e-11    2
-.271428065e+06-.474657811e+04-.269350780e+03 .391998234e+01-.105525918e-02    3
-.168858987e-05 .972637936e-09 .722971705e+05 .141824356e+04                   4
BIN6C                   C 640H  34          G   300.00   4000.00  1000.00      1
 .816745766e+03 .130541967e+01-.482467007e-03 .803609911e-07-.499915059e-11    2
-.420769482e+06-.454055202e+04-.260894565e+03 .353895191e+01-.666844909e-03    3
-.190047075e-05 .100428001e-08-.105083869e+06 .117013783e+04                   4
BIN7A                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          813
 .227996401e+04 .364410804e+01-.134681737e-02 .224329490e-06-.139552395e-10    2
 .219703936e+06-.125294003e+05-.798183644e+03 .125608657e+02-.983885162e-02    3
 .263510017e-05 .228737231e-09 .101891965e+07 .319868647e+04                   4
BIN7B                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          250
 .174821343e+04 .279420142e+01-.103270238e-02 .172009660e-06-.107004925e-10    2
-.528501603e+06-.927449889e+04-.525643684e+03 .765707323e+01-.206469049e-02    3
-.329407582e-05 .189828623e-08 .142639667e+06 .276398698e+04                   4
BIN7C                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H           65
 .159398623e+04 .254769728e+01-.941597491e-03 .156834989e-06-.975649647e-11    2
-.824746508e+06-.886326423e+04-.509649220e+03 .690588633e+01-.129480205e-02    3
-.371700233e-05 .196265639e-08-.208493980e+06 .228472375e+04                   4
BIN8A                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H         1563
 .452144611e+04 .722670975e+01-.267090277e-02 .444872681e-06-.276749385e-10    2
 .525439399e+06-.253601694e+05-.163861142e+04 .254934056e+02-.207827201e-01    3
 .632122666e-05 .101241844e-09 .209454960e+07 .599019956e+04                   4
BIN8B                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          500
 .349623033e+04 .558808872e+01-.206528866e-02 .343999983e-06-.213997822e-10    2
-.106037670e+07-.185413207e+05-.105215148e+04 .153124310e+02-.412210619e-02    3
-.659605418e-05 .379936694e-08 .282300003e+06 .554001391e+04                   4
BIN8C                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          126
 .318473927e+04 .509022690e+01-.188128508e-02 .313351859e-06-.194932032e-10    2
-.165413482e+07-.177215999e+05-.101850654e+04 .137964163e+02-.257671322e-02    3
-.743906960e-05 .392526201e-08-.423020017e+06 .455286982e+04                   4
BIN9A                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         3000
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .105415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .433609933e+07 .163588732e+05                   4
BIN9B                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         1000
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.212075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .564600007e+06 .110800278e+05                   4
BIN9C                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          251
 .636869480e+04 .101792011e+02-.376210719e-02 .626626605e-06-.389816093e-10    2
-.330896407e+07-.354429274e+05-.203670710e+04 .275892080e+02-.515111307e-02    3
-.148784176e-04 .785016202e-08-.847131304e+06 .910009023e+04                   4
BIN10A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5750
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .171313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .820225091e+07 .320518708e+05                   4
BIN10B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         2000
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.424150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .112920001e+07 .221600556e+05                   4
BIN10C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          501
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.662199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.169833321e+07 .182065710e+05                   4
BIN11A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        11000
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .262917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .154586477e+08 .627960702e+05                   4
BIN11B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         4000
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.848301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .225840003e+07 .443201113e+05                   4
BIN11C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1001
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.132446866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.339775769e+07 .364074926e+05                   4
BIN12A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        21000
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .367089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290315457e+08 .122952718e+06                   4
BIN12B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         8000
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169660271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .451680005e+07 .886402226e+05                   4
BIN12C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2001
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264900676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.679660664e+07 .728093358e+05                   4
BIN13A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        40000
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .416688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .542915920e+08 .240626590e+06                   4
BIN13B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        16000
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.339320543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .903360011e+07 .177280445e+06                   4
BIN13C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4001
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529808296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135943046e+08 .145613022e+06                   4
BIN14A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        76000
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .198394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101040185e+09 .470695489e+06                   4
BIN14B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        32000
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678641086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .180672002e+08 .354560890e+06                   4
BIN14C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8001
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105962354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271897004e+08 .291220395e+06                   4
BIN15A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       144000
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.873175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .186994373e+09 .920275597e+06                   4
BIN15B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        64000
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135728217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361344004e+08 .709121781e+06                   4
BIN15C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16001
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211925402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543804920e+08 .582435141e+06                   4
BIN16A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       272000
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428627973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343816752e+09 .179832043e+07                   4
BIN16B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       128000
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271456434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .722688009e+08 .141824356e+07                   4
BIN16C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32001
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423851498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108762075e+09 .116486463e+07                   4
BIN17A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       500000
 .195633111e+07 .312683969e+04-.115564137e+01 .192486706e-03-.119743423e-07    2
-.133324395e+09-.981860207e+07-.548565677e+06 .866959432e+04-.309406979e+01    3
-.273451411e-02 .181552901e-05 .612587417e+09 .342986263e+07                   4
BIN17B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       250000
 .174811516e+07 .279404436e+04-.103264433e+01 .171999992e-03-.106998911e-07    2
-.530188348e+09-.927066036e+07-.526075742e+06 .765621551e+04-.206105310e+01    3
-.329802709e-02 .189968347e-05 .141150002e+09 .277000696e+07                   4
BIN17C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H        62501
 .159195398e+07 .254444911e+04-.940397008e+00 .156635033e-03-.974405749e-08    2
-.827835618e+09-.885970435e+07-.509208597e+06 .689618503e+04-.128629289e+01    3
-.372066155e-02 .196279968e-05-.212426969e+09 .227512085e+07                   4
BIN18A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       937500
 .386060824e+07 .617048055e+04-.228053348e+01 .379851734e-03-.236300717e-07    2
-.365864779e+09-.195002187e+08-.109150887e+07 .170858439e+05-.592988540e+01    3
-.560990646e-02 .365209663e-05 .110731548e+10 .669476134e+07                   4
BIN18B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       500000
 .349623033e+07 .558808872e+04-.206528866e+01 .343999983e-03-.213997822e-07    2
-.106037670e+10-.185413207e+08-.105215148e+07 .153124310e+05-.412210619e+01    3
-.659605418e-02 .379936694e-05 .282300003e+09 .554001391e+07                   4
BIN18C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       125001
 .318390719e+07 .508889697e+04-.188079355e+01 .313269989e-03-.194881102e-07    2
-.165567193e+10-.177194084e+08-.101841689e+07 .137923664e+05-.257258347e+01    3
-.744132337e-02 .392559899e-05-.424855028e+09 .455023605e+07                   4
BIN19A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H      1750000
 .761710851e+07 .121745634e+05-.449956845e+01 .749460110e-03-.466229179e-07    2
-.930161534e+09-.387264666e+08-.217177277e+07 .336649985e+05-.113432625e+02    3
-.115015694e-01 .734627050e-05 .197891225e+10 .130595948e+08                   4
BIN19B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H      1000000
 .699246065e+07 .111761774e+05-.413057731e+01 .687999967e-03-.427995643e-07    2
-.212075339e+10-.370826415e+08-.210430297e+07 .306248620e+05-.824421238e+01    3
-.131921084e-01 .759873388e-05 .564600007e+09 .110800278e+08                   4
BIN19C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H       250001
 .636781359e+07 .101777927e+05-.376158664e+01 .626539901e-03-.389762156e-07    2
-.331134456e+10-.354388166e+08-.203683347e+07 .275847292e+05-.514516462e+01    3
-.148826470e-01 .785119762e-05-.849711148e+09 .910046645e+07                   4
BIN20A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      3250000
 .150260011e+08 .240163315e+05-.887613985e+01 .147843351e-02-.919713846e-07    2
-.225718702e+10-.769049915e+08-.432105561e+07 .663166181e+05-.216535082e+02    3
-.235666518e-01 .147766955e-04 .348638709e+10 .254593340e+08                   4
BIN20B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      2000000
 .139849213e+08 .223523549e+05-.826115463e+01 .137599993e-02-.855991287e-07    2
-.424150678e+10-.741652829e+08-.420860594e+07 .612497241e+05-.164884248e+02    3
-.263842167e-01 .151974678e-04 .112920001e+10 .221600556e+08                   4
BIN20C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H       500001
 .127356264e+08 .203555841e+05-.752317282e+01 .125307972e-02-.779524263e-07    2
-.662268981e+10-.708776329e+08-.407366664e+07 .551694548e+05-.102903269e+02    3
-.297652943e-01 .157023949e-04-.169942339e+10 .182009272e+08                   4
BIN21A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      6000000
 .296355702e+08 .473670724e+05-.175062856e+02 .291589358e-02-.181393867e-06    2
-.530810195e+10-.152714099e+09-.859713135e+07 .130606479e+06-.412409831e+02    3
-.482603296e-01 .297216998e-04 .602989935e+10 .495989567e+08                   4
BIN21B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      4000000
 .279698426e+08 .447047097e+05-.165223093e+02 .275199987e-02-.171198257e-06    2
-.848301357e+10-.148330566e+09-.841721188e+07 .122499448e+06-.329768495e+02    3
-.527684334e-01 .303949355e-04 .225840003e+10 .443201113e+08                   4
BIN21C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      1000001
 .254712520e+08 .407111670e+05-.150463452e+02 .250615937e-02-.155904848e-06    2
-.132453803e+11-.141755266e+09-.814733297e+07 .110338906e+06-.205806515e+02    3
-.595305889e-01 .314047894e-04-.339884787e+10 .364018488e+08                   4
BIN22A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H     12000000
 .592711404e+08 .947341447e+05-.350125712e+02 .583178717e-02-.362787734e-06    2
-.106162039e+11-.305428199e+09-.171942627e+08 .261212957e+06-.824819661e+02    3
-.965206591e-01 .594433996e-04 .120597987e+11 .991979134e+08                   4
BIN22B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      8000000
 .559396852e+08 .894094194e+05-.330446185e+02 .550399973e-02-.342396515e-06    2
-.169660271e+11-.296661132e+09-.168344238e+08 .244998896e+06-.659536990e+02    3
-.105536867e+00 .607898710e-04 .451680005e+10 .886402226e+08                   4
BIN22C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      2000001
 .509425024e+08 .814223315e+05-.300926894e+02 .501231859e-02-.311809686e-06    2
-.264907620e+11-.283510531e+09-.162946653e+08 .220677805e+06-.411612984e+02    3
-.119061178e+00 .628095780e-04-.679769791e+10 .728036864e+08                   4
BIN23A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     24000000
 .118542281e+09 .189468289e+06-.700251424e+02 .116635743e-01-.725575467e-06    2
-.212324078e+11-.610856398e+09-.343885254e+08 .522425915e+06-.164963932e+03    3
-.193041318e+00 .118886799e-03 .241195974e+11 .198395827e+09                   4
BIN23B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     16000000
 .111879370e+09 .178818839e+06-.660892370e+02 .110079995e-01-.684793029e-06    2
-.339320543e+11-.593322263e+09-.336688475e+08 .489997793e+06-.131907398e+03    3
-.211073734e+00 .121579742e-03 .903360011e+10 .177280445e+09                   4
BIN23C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H      4000001
 .101885006e+09 .162844664e+06-.601853793e+02 .100246373e-01-.623619377e-06    2
-.529815233e+11-.567021061e+09-.325893310e+08 .441355613e+06-.823225992e+02    3
-.238122356e+00 .125619156e-03-.135953947e+11 .145607378e+09                   4
BIN24A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     48000000
 .237084562e+09 .378936579e+06-.140050285e+03 .233271487e-01-.145115093e-05    2
-.424648156e+11-.122171280e+10-.687770508e+08 .104485183e+07-.329927864e+03    3
-.386082637e+00 .237773599e-03 .482391948e+11 .396791654e+09                   4
BIN24B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     32000000
 .223758741e+09 .357637678e+06-.132178474e+03 .220159989e-01-.136958606e-05    2
-.678641086e+11-.118664453e+10-.673376950e+08 .979995585e+06-.263814796e+03    3
-.422147467e+00 .243159484e-03 .180672002e+11 .354560890e+09                   4
BIN24C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H      8000001
 .203770010e+09 .325689327e+06-.120370758e+03 .200492744e-01-.124723875e-05    2
-.105963047e+12-.113404212e+10-.651786616e+08 .882711223e+06-.164645196e+03    3
-.476244713e+00 .251238313e-03-.271907906e+11 .291214751e+09                   4
BIN25A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     96000000
 .474169124e+09 .757873158e+06-.280100570e+03 .466542973e-01-.290230187e-05    2
-.849296311e+11-.244342559e+10-.137554102e+09 .208970366e+07-.659855729e+03    3
-.772165273e+00 .475547197e-03 .964783896e+11 .793583307e+09                   4
BIN25B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     64000000
 .447517482e+09 .715275356e+06-.264356948e+03 .440319979e-01-.273917212e-05    2
-.135728217e+12-.237328905e+10-.134675390e+09 .195999117e+07-.527629592e+03    3
-.844294935e+00 .486318968e-03 .361344004e+11 .709121781e+09                   4
BIN25C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     16000001
 .407540020e+09 .651378653e+06-.240741516e+03 .400985488e-01-.249447749e-05    2
-.211926095e+12-.226808425e+10-.130357323e+09 .176542244e+07-.329290390e+03    3
-.952489427e+00 .502476625e-03-.543815822e+11 .582429497e+09                   4
BIN1AJ                  C  20H  15          G   300.00   4000.00  1000.00      1
 .384004130e+02 .613760802e-01-.226838420e-04 .377828116e-08-.235041851e-12    2
 .583425289e+05-.190858878e+03-.946290891e+01 .179252381e+00-.989756752e-04    3
-.116559979e-07 .214782048e-10 .722142317e+05 .597553003e+02                   4
BIN1BJ                  C  20H   9          G   300.00   4000.00  1000.00      1
 .329670254e+02 .526917977e-01-.194742383e-04 .324368101e-08-.201785086e-12    2
 .610771833e+05-.161481167e+03-.895697031e+01 .146820540e+00-.577692501e-04    3
-.392441219e-07 .283752285e-10 .736083600e+05 .601566475e+02                   4
BIN1CJ                  C  20H   4          G   300.00   4000.00  1000.00      1
 .288518394e+02 .461144212e-01-.170433212e-04 .283878100e-08-.176596796e-12    2
 .538768910e+05-.152441597e+03-.829114243e+01 .126981825e+00-.389276128e-04    3
-.485387475e-07 .293596977e-10 .648180581e+05 .439495435e+02                   4
BIN2AJ                  C  40H  30          G   300.00   4000.00  1000.00      1
 .759883346e+02 .121453540e+00-.448877300e-04 .747661988e-08-.465110589e-12    2
 .603973953e+05-.376351286e+03-.224069955e+02 .373191638e+00-.228373343e-03    3
 .179614865e-08 .353583380e-10 .883409758e+05 .136281912e+03                   4
BIN2BJ                  C  40H  15          G   300.00   4000.00  1000.00      1
 .626025956e+02 .100058870e+00-.369805239e-04 .615957460e-08-.383178953e-12    2
 .556485106e+05-.314195266e+03-.175541017e+02 .277427018e+00-.990102332e-04    3
-.875044514e-07 .580969283e-10 .795176885e+05 .109755604e+03                   4
BIN2CJ                  C  40H   7          G   300.00   4000.00  1000.00      1
 .559396852e+02 .894094194e-01-.330446185e-04 .550399973e-08-.342396515e-12    2
 .429914185e+05-.296661132e+03-.168344238e+02 .244998896e+00-.659536990e-04    3
-.105536867e-06 .607898710e-10 .644742457e+05 .886402226e+02                   4
BIN3AJ                  C  80H  59          G   300.00   4000.00  1000.00      1
 .150797478e+03 .241022357e+00-.890788896e-04 .148372172e-07-.923003567e-12    2
 .630318960e+05-.764406699e+03-.455633619e+02 .756332498e+00-.489114578e-03    3
 .351844886e-07 .598168799e-10 .117848100e+06 .254746237e+03                   4
BIN3BJ                  C  80H  23          G   300.00   4000.00  1000.00      1
 .118542281e+03 .189468289e+00-.700251424e-04 .116635743e-07-.725575467e-12    2
 .386399290e+05-.610856398e+03-.343885254e+02 .522425915e+00-.164963932e-03    3
-.193041318e-06 .118886799e-09 .839919342e+05 .198395827e+03                   4
BIN3CJ                  C  80H   7          G   300.00   4000.00  1000.00      1
 .105216460e+03 .168169388e+00-.621533316e-04 .103524246e-07-.644010591e-12    2
 .133257448e+05-.575788129e+03-.329491696e+02 .457569671e+00-.988508639e-04    3
-.229106149e-06 .124272685e-09 .539050484e+05 .156165064e+03                   4
BIN4AJ                  C 160H 115          G   300.00   4000.00  1000.00      1
 .299236573e+03 .478275269e+00-.176764639e-03 .294423892e-07-.183157191e-11    2
 .705380025e+05-.155222165e+04-.926254655e+02 .153256344e+01-.104296494e-02    3
 .133553360e-06 .978341677e-10 .178028497e+06 .473857298e+03                   4
BIN4BJ                  C 160H  31          G   300.00   4000.00  1000.00      1
 .223758741e+03 .357637678e+00-.132178474e-03 .220159989e-07-.136958606e-11    2
-.803432616e+04-.118664453e+04-.673376950e+02 .979995585e+00-.263814796e-03    3
-.422147467e-06 .243159484e-09 .778969826e+05 .354560890e+03                   4
BIN4CJ                  C 160H   9          G   300.00   4000.00  1000.00      1
 .205435737e+03 .328351689e+00-.121354734e-03 .202131681e-07-.125743435e-11    2
-.427526744e+05-.113842566e+04-.653585808e+02 .890818250e+00-.172909327e-03    3
-.471736610e-06 .250565077e-09 .366161697e+05 .296493591e+03                   4
BIN5AJ                  C 320H 223          G   300.00   4000.00  1000.00      1
 .593310588e+03 .948299129e+00-.350479658e-03 .583768256e-07-.363154476e-11    2
 .952119959e+05-.312882274e+04-.194461399e+03 .312434830e+01-.224387754e-02    3
 .412099583e-06 .147772804e-09 .307380465e+06 .927804457e+03                   4
BIN5BJ                  C 320H  63          G   300.00   4000.00  1000.00      1
 .447517482e+03 .715275356e+00-.264356948e-03 .440319979e-07-.273917212e-11    2
-.757140323e+05-.237328905e+04-.134675390e+03 .195999117e+01-.527629592e-03    3
-.844294935e-06 .486318968e-09 .961485852e+05 .709121781e+03                   4
BIN5CJ                  C 320H  17          G   300.00   4000.00  1000.00      1
 .409205747e+03 .654041015e+00-.241725492e-03 .402624424e-07-.250467310e-11    2
-.148758277e+06-.227246778e+04-.130537242e+03 .177352947e+01-.337554521e-03    3
-.947981323e-06 .501803389e-09 .938282361e+04 .587708337e+03                   4
BIN6AJ                  C 640H 431          G   300.00   4000.00  1000.00      1
 .117696475e+04 .188116422e+01-.695255086e-03 .115803539e-06-.720398434e-11    2
 .150914619e+06-.634005997e+04-.398024258e+03 .633800264e+01-.476093625e-02    3
 .108624875e-05 .206199066e-09 .567419557e+06 .173874832e+04                   4
BIN6BJ                  C 640H 127          G   300.00   4000.00  1000.00      1
 .895034964e+03 .143055071e+01-.528713896e-03 .880639958e-07-.547834423e-11    2
-.211428065e+06-.474657811e+04-.269350780e+03 .391998234e+01-.105525918e-02    3
-.168858987e-05 .972637936e-09 .132297170e+06 .141824356e+04                   4
BIN6CJ                  C 640H  33          G   300.00   4000.00  1000.00      1
 .816745766e+03 .130541967e+01-.482467007e-03 .803609911e-07-.499915059e-11    2
-.360769482e+06-.454055202e+04-.260894565e+03 .353895191e+01-.666844909e-03    3
-.190047075e-05 .100428001e-08-.450838685e+05 .117013783e+04                   4
BIN7AJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          812
 .227996401e+04 .364410804e+01-.134681737e-02 .224329490e-06-.139552395e-10    2
 .279703936e+06-.125294003e+05-.798183644e+03 .125608657e+02-.983885162e-02    3
 .263510017e-05 .228737231e-09 .107891965e+07 .319868647e+04                   4
BIN7BJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          249
 .174821343e+04 .279420142e+01-.103270238e-02 .172009660e-06-.107004925e-10    2
-.468501603e+06-.927449889e+04-.525643684e+03 .765707323e+01-.206469049e-02    3
-.329407582e-05 .189828623e-08 .202639667e+06 .276398698e+04                   4
BIN7CJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H           64
 .159398623e+04 .254769728e+01-.941597491e-03 .156834989e-06-.975649647e-11    2
-.764746508e+06-.886326423e+04-.509649220e+03 .690588633e+01-.129480205e-02    3
-.371700233e-05 .196265639e-08-.148493980e+06 .228472375e+04                   4
BIN8AJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H         1562
 .452144611e+04 .722670975e+01-.267090277e-02 .444872681e-06-.276749385e-10    2
 .585439399e+06-.253601694e+05-.163861142e+04 .254934056e+02-.207827201e-01    3
 .632122666e-05 .101241844e-09 .215454960e+07 .599019956e+04                   4
BIN8BJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          499
 .349623033e+04 .558808872e+01-.206528866e-02 .343999983e-06-.213997822e-10    2
-.100037670e+07-.185413207e+05-.105215148e+04 .153124310e+02-.412210619e-02    3
-.659605418e-05 .379936694e-08 .342300003e+06 .554001391e+04                   4
BIN8CJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          125
 .318473927e+04 .509022690e+01-.188128508e-02 .313351859e-06-.194932032e-10    2
-.159413482e+07-.177215999e+05-.101850654e+04 .137964163e+02-.257671322e-02    3
-.743906960e-05 .392526201e-08-.363020017e+06 .455286982e+04                   4
BIN9AJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         2999
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .111415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .439609933e+07 .163588732e+05                   4
BIN9BJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          999
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.206075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .624600007e+06 .110800278e+05                   4
BIN9CJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          250
 .636869480e+04 .101792011e+02-.376210719e-02 .626626605e-06-.389816093e-10    2
-.324896407e+07-.354429274e+05-.203670710e+04 .275892080e+02-.515111307e-02    3
-.148784176e-04 .785016202e-08-.787131304e+06 .910009023e+04                   4
BIN10AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5749
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .177313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .826225091e+07 .320518708e+05                   4
BIN10BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         1999
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.418150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .118920001e+07 .221600556e+05                   4
BIN10CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          500
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.656199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.163833321e+07 .182065710e+05                   4
BIN11AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        10999
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .268917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .155186477e+08 .627960702e+05                   4
BIN11BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         3999
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.842301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .231840003e+07 .443201113e+05                   4
BIN11CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1000
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.131846866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.333775769e+07 .364074926e+05                   4
BIN12AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        20999
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .373089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290915457e+08 .122952718e+06                   4
BIN12BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         7999
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169060271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .457680005e+07 .886402226e+05                   4
BIN12CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2000
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264300676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.673660664e+07 .728093358e+05                   4
BIN13AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        39999
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .422688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .543515920e+08 .240626590e+06                   4
BIN13BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        15999
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.338720543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .909360011e+07 .177280445e+06                   4
BIN13CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4000
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529208296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135343046e+08 .145613022e+06                   4
BIN14AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        75999
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .204394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101100185e+09 .470695489e+06                   4
BIN14BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        31999
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678041086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .181272002e+08 .354560890e+06                   4
BIN14CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8000
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105902354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271297004e+08 .291220395e+06                   4
BIN15AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       143999
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.867175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .187054373e+09 .920275597e+06                   4
BIN15BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        63999
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135668217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361944004e+08 .709121781e+06                   4
BIN15CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16000
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211865402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543204920e+08 .582435141e+06                   4
BIN16AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       271999
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428027973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343876752e+09 .179832043e+07                   4
BIN16BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       127999
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271396434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .723288009e+08 .141824356e+07                   4
BIN16CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32000
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423791498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108702075e+09 .116486463e+07                   4
BIN17AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       499999
 .195633111e+07 .312683969e+04-.115564137e+01 .192486706e-03-.119743423e-07    2
-.133264395e+09-.981860207e+07-.548565677e+06 .866959432e+04-.309406979e+01    3
-.273451411e-02 .181552901e-05 .612647417e+09 .342986263e+07                   4
BIN17BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       249999
 .174811516e+07 .279404436e+04-.103264433e+01 .171999992e-03-.106998911e-07    2
-.530128348e+09-.927066036e+07-.526075742e+06 .765621551e+04-.206105310e+01    3
-.329802709e-02 .189968347e-05 .141210002e+09 .277000696e+07                   4
BIN17CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H        62500
 .159195398e+07 .254444911e+04-.940397008e+00 .156635033e-03-.974405749e-08    2
-.827775618e+09-.885970435e+07-.509208597e+06 .689618503e+04-.128629289e+01    3
-.372066155e-02 .196279968e-05-.212366969e+09 .227512085e+07                   4
BIN18AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       937499
 .386060824e+07 .617048055e+04-.228053348e+01 .379851734e-03-.236300717e-07    2
-.365804779e+09-.195002187e+08-.109150887e+07 .170858439e+05-.592988540e+01    3
-.560990646e-02 .365209663e-05 .110737548e+10 .669476134e+07                   4
BIN18BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       499999
 .349623033e+07 .558808872e+04-.206528866e+01 .343999983e-03-.213997822e-07    2
-.106031670e+10-.185413207e+08-.105215148e+07 .153124310e+05-.412210619e+01    3
-.659605418e-02 .379936694e-05 .282360003e+09 .554001391e+07                   4
BIN18CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       125000
 .318390719e+07 .508889697e+04-.188079355e+01 .313269989e-03-.194881102e-07    2
-.165561193e+10-.177194084e+08-.101841689e+07 .137923664e+05-.257258347e+01    3
-.744132337e-02 .392559899e-05-.424795028e+09 .455023605e+07                   4
BIN19AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H      1749999
 .761710851e+07 .121745634e+05-.449956845e+01 .749460110e-03-.466229179e-07    2
-.930101534e+09-.387264666e+08-.217177277e+07 .336649985e+05-.113432625e+02    3
-.115015694e-01 .734627050e-05 .197897225e+10 .130595948e+08                   4
BIN19BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H       999999
 .699246065e+07 .111761774e+05-.413057731e+01 .687999967e-03-.427995643e-07    2
-.212069339e+10-.370826415e+08-.210430297e+07 .306248620e+05-.824421238e+01    3
-.131921084e-01 .759873388e-05 .564660007e+09 .110800278e+08                   4
BIN19CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H       250000
 .636781359e+07 .101777927e+05-.376158664e+01 .626539901e-03-.389762156e-07    2
-.331128456e+10-.354388166e+08-.203683347e+07 .275847292e+05-.514516462e+01    3
-.148826470e-01 .785119762e-05-.849651148e+09 .910046645e+07                   4
BIN20AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      3249999
 .150260011e+08 .240163315e+05-.887613985e+01 .147843351e-02-.919713846e-07    2
-.225712702e+10-.769049915e+08-.432105561e+07 .663166181e+05-.216535082e+02    3
-.235666518e-01 .147766955e-04 .348644709e+10 .254593340e+08                   4
BIN20BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      1999999
 .139849213e+08 .223523549e+05-.826115463e+01 .137599993e-02-.855991287e-07    2
-.424144678e+10-.741652829e+08-.420860594e+07 .612497241e+05-.164884248e+02    3
-.263842167e-01 .151974678e-04 .112926001e+10 .221600556e+08                   4
BIN20CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H       500000
 .127356264e+08 .203555841e+05-.752317282e+01 .125307972e-02-.779524263e-07    2
-.662262981e+10-.708776329e+08-.407366664e+07 .551694548e+05-.102903269e+02    3
-.297652943e-01 .157023949e-04-.169936339e+10 .182009272e+08                   4
BIN21AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      5999999
 .296355702e+08 .473670724e+05-.175062856e+02 .291589358e-02-.181393867e-06    2
-.530804195e+10-.152714099e+09-.859713135e+07 .130606479e+06-.412409831e+02    3
-.482603296e-01 .297216998e-04 .602995935e+10 .495989567e+08                   4
BIN21BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      3999999
 .279698426e+08 .447047097e+05-.165223093e+02 .275199987e-02-.171198257e-06    2
-.848295357e+10-.148330566e+09-.841721188e+07 .122499448e+06-.329768495e+02    3
-.527684334e-01 .303949355e-04 .225846003e+10 .443201113e+08                   4
BIN21CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      1000000
 .254712520e+08 .407111670e+05-.150463452e+02 .250615937e-02-.155904848e-06    2
-.132453203e+11-.141755266e+09-.814733297e+07 .110338906e+06-.205806515e+02    3
-.595305889e-01 .314047894e-04-.339878787e+10 .364018488e+08                   4
BIN22AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H     11999999
 .592711404e+08 .947341447e+05-.350125712e+02 .583178717e-02-.362787734e-06    2
-.106161439e+11-.305428199e+09-.171942627e+08 .261212957e+06-.824819661e+02    3
-.965206591e-01 .594433996e-04 .120598587e+11 .991979134e+08                   4
BIN22BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      7999999
 .559396852e+08 .894094194e+05-.330446185e+02 .550399973e-02-.342396515e-06    2
-.169659671e+11-.296661132e+09-.168344238e+08 .244998896e+06-.659536990e+02    3
-.105536867e+00 .607898710e-04 .451686005e+10 .886402226e+08                   4
BIN22CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      2000000
 .509425024e+08 .814223315e+05-.300926894e+02 .501231859e-02-.311809686e-06    2
-.264907020e+11-.283510531e+09-.162946653e+08 .220677805e+06-.411612984e+02    3
-.119061178e+00 .628095780e-04-.679763791e+10 .728036864e+08                   4
BIN23AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     23999999
 .118542281e+09 .189468289e+06-.700251424e+02 .116635743e-01-.725575467e-06    2
-.212323478e+11-.610856398e+09-.343885254e+08 .522425915e+06-.164963932e+03    3
-.193041318e+00 .118886799e-03 .241196574e+11 .198395827e+09                   4
BIN23BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     15999999
 .111879370e+09 .178818839e+06-.660892370e+02 .110079995e-01-.684793029e-06    2
-.339319943e+11-.593322263e+09-.336688475e+08 .489997793e+06-.131907398e+03    3
-.211073734e+00 .121579742e-03 .903366011e+10 .177280445e+09                   4
BIN23CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H      4000000
 .101885006e+09 .162844664e+06-.601853793e+02 .100246373e-01-.623619377e-06    2
-.529814633e+11-.567021061e+09-.325893310e+08 .441355613e+06-.823225992e+02    3
-.238122356e+00 .125619156e-03-.135953347e+11 .145607378e+09                   4
BIN24AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     47999999
 .237084562e+09 .378936579e+06-.140050285e+03 .233271487e-01-.145115093e-05    2
-.424647556e+11-.122171280e+10-.687770508e+08 .104485183e+07-.329927864e+03    3
-.386082637e+00 .237773599e-03 .482392548e+11 .396791654e+09                   4
BIN24BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     31999999
 .223758741e+09 .357637678e+06-.132178474e+03 .220159989e-01-.136958606e-05    2
-.678640486e+11-.118664453e+10-.673376950e+08 .979995585e+06-.263814796e+03    3
-.422147467e+00 .243159484e-03 .180672602e+11 .354560890e+09                   4
BIN24CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H      8000000
 .203770010e+09 .325689327e+06-.120370758e+03 .200492744e-01-.124723875e-05    2
-.105962987e+12-.113404212e+10-.651786616e+08 .882711223e+06-.164645196e+03    3
-.476244713e+00 .251238313e-03-.271907306e+11 .291214751e+09                   4
BIN25AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     95999999
 .474169124e+09 .757873158e+06-.280100570e+03 .466542973e-01-.290230187e-05    2
-.849295711e+11-.244342559e+10-.137554102e+09 .208970366e+07-.659855729e+03    3
-.772165273e+00 .475547197e-03 .964784496e+11 .793583307e+09                   4
BIN25BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     63999999
 .447517482e+09 .715275356e+06-.264356948e+03 .440319979e-01-.273917212e-05    2
-.135728157e+12-.237328905e+10-.134675390e+09 .195999117e+07-.527629592e+03    3
-.844294935e+00 .486318968e-03 .361344604e+11 .709121781e+09                   4
BIN25CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     16000000
 .407540020e+09 .651378653e+06-.240741516e+03 .400985488e-01-.249447749e-05    2
-.211926035e+12-.226808425e+10-.130357323e+09 .176542244e+07-.329290390e+03    3
-.952489427e+00 .502476625e-03-.543815222e+11 .582429497e+09                   4
! Kik add C6H4C2H3 radical from Burcat A1C2H3*
C6H4C2H3          T12/07C  8.H  7.   0.   0.G   200.000  6000.000 1000.00      1
 1.57334515E+01 2.38965492E-02-8.60829763E-06 1.39223384E-09-8.35065775E-14    2
 4.08827573E+04-5.82476667E+01 1.17830774E+00 3.40765502E-02 5.85065530E-05    3
-1.10953244E-07 4.95222636E-11 4.61414992E+04 2.36053284E+01 4.83284254E+04    4
!Blanq A1C2H3Y
!C6H4C2H3          000000N   0H   7O   0C   8G       300      3000    1000      1
! 3.90114779E+00 5.15894020E-02-3.05080522E-05 8.55910896E-09-9.23046757E-13    2
! 4.59935428E+04 5.96930655E+00-5.36214520E+00 8.67033297E-02-7.54297960E-05    3
! 3.01139854E-08-3.40681418E-12 4.77818209E+04 5.07407949E+01                   4
!KAUST
!A1C2H3*           000000N   0H   7O   0C   8G       300      3000    1000      1
! 3.90114779E+00 5.15894020E-02-3.05080522E-05 8.55910896E-09-9.23046757E-13    2
! 4.59935428E+04 5.96930655E+00-5.36214520E+00 8.67033297E-02-7.54297960E-05    3
! 3.01139854E-08-3.40681418E-12 4.77818209E+04 5.07407949E+01                   4
!
! Add all intermediates from burcat
!1-naphthyl-W2           C  10H   7          G    300.00   4000.00 1000.00      1
! .146529084E+02 .356159360E-01-.121796480E-04 .138747960E-08 .000000000E+00    2
! .405898415E+05-.575649187E+02-.631700500E+01 .913910790E-01-.608201990E-04    3
! .152228010E-07 .000000000E+00 .464268700E+05 .512234700E+02                   4
!2-naphthyl-W4           C  10H   7          G    300.00   4000.00 1000.00      1
! .146529084E+02 .356159360E-01-.121796480E-04 .138747960E-08 .000000000E+00    2
! .405898415E+05-.575649187E+02-.631700500E+01 .913910790E-01-.608201990E-04    3
! .152228010E-07 .000000000E+00 .464268700E+05 .512234700E+02                   4
!RA1R5CH3
!
!
!
naphthyne12       T 7/98C 10.H  6.   0.   0.G   200.000  6000.000 3000.0       1
 1.87728941E+01 2.48768793E-02-9.09940935E-06 1.48730676E-09-8.98228135E-14    2
 5.15727443E+04-7.68608875E+01-1.50617131E+00 6.03325879E-02 1.09063952E-05    3
-6.91994009E-08 3.54144371E-11 5.80261788E+04 3.24494940E+01 6.02350349E+04    4
naphthyne23       T 7/98C 10.H  6.   0.   0.G   200.000  6000.000 3000.0       1
 1.87728941E+01 2.48768793E-02-9.09940935E-06 1.48730676E-09-8.98228135E-14    2
 5.15727443E+04-7.68608875E+01-1.50617131E+00 6.03325879E-02 1.09063952E-05    3
-6.91994009E-08 3.54144371E-11 5.80261788E+04 3.24494940E+01 6.02350349E+04    4
!
!126738-27-0 or 182180-84-3
!C10H9 phenyl-butadienyl radical C6H5-CH=CH-CH=CH*  SIGMA=1  STATWT=2  IA=17.2514
!IB=140.1877  IC=157.4391  Ir(-CH=CH-CH=CH*)=7.03118  ROSYM=1  V(3)=1224. cm-1
!est.  Ir(-CH=CH*)=2.59427  ROSYM=1  V(3)524. cm-1 as in butadiene.  Nu=3268,
!3212,3204,3195,3186,3183,3176,3144,3040,1693,1661,1645,1631,1546,1497,1380,1372,
!1343,1321,1253,1249,1218,1193,1162,1112,1060,1015,1013,991,964,927,889,859,852,
!832(2),768,705,639,635,621,513,510,414,343,313,297,174.8,124.54   HF298=106.24
!kcal  REF=Thergas   c(#1)&ch&ch&ch&ch&ch&1,1/ch//ch//ch//ch(.)   {HF298=106.5
!kcal  REF=NIST 94}  Max Lst Sq Error Cp @ 200 K 0.66%
C6H5CHCHCHCH         /06C 10.H  9.   0.   0.G   200.000  6000.000 3000.0       1 
 1.97227364E+01 3.05121625E-02-1.10537483E-05 1.79050874E-09-1.07387763E-13    2
 4.42281159E+04-7.53736816E+01 2.29508183E+00 4.52323197E-02 5.98076375E-05    3
-1.21133405E-07 5.46626377E-11 5.04522033E+04 2.21435730E+01 5.34617386E+04    4
!1785-61-1
!C10H6 1,3-diethynylBenzene 1,3-C6H4(CCH)2  SIGMA=2  STATWT=1  IA=31.252
!IB=92.9373  IC=124.1894  Nu=115,126,162,186,368,388,465,469,500,505,561,572,576,
!629.5(2),646,702,718,812,916,921,925,983,1014,1122,1175,1205,1273,1313.5,1355,
!1446,1525,1623,1649,2227.6(2),3197,3216,3223,3228,3494.3(2)  HF298=131.96+/-2.
!kcal  REF=Elke Goos G3B3  Max Lst Sq Error Cp @ 1300 K 0.47%.
C6H4(C2H)2        T10/15C 10.H  6.   0.   0.G   200.000  6000.000 3000.0       1
 1.94890277E+01 2.35101034E-02-8.43787249E-06 1.36207463E-09-8.15578305E-14    2
 5.80245053E+04-7.66298995E+01-1.92263481E+00 8.57578670E-02-7.03095425E-05    3
 2.10427011E-08 1.27338464E-12 6.37450309E+04 3.30657524E+01 6.64044712E+04    4
! Fei Qi
! Benzofulvene
!C9H6CH2   MATSUGI2013   C  10H   8    0    0G   300.000  5000.000 1401.00      1
Benzofulvene            C  10H   8    0    0G   300.000  5000.000 1401.00      1
 2.37888939E+01 2.39146033E-02-8.24877665E-06 1.28829948E-09-7.50678039E-14    2
 1.43968777E+04-1.07094280E+02-8.01337918E+00 1.08401947E-01-9.55671696E-05    3
 4.25996671E-08-7.54462202E-12 2.43488603E+04 5.99659944E+01                   4
!benzofulvenyl radical
!C9H7CH2   MATSUGI2013   C  10H   9    0    0G   300.000  5000.000 1400.00      1
! 2.48973930E+01 2.55147986E-02-8.79922194E-06 1.37404921E-09-8.00535169E-14    2
! 1.83072953E+04-1.12654689E+02-8.02975915E+00 1.12889393E-01-9.91274443E-05    3
! 4.41732177E-08-7.83596047E-12 2.86367245E+04 6.03761192E+01                   4
!536738-49-5
!C10H9 1-methyl-1-indenyl Radical  SIGMA=1 STATWT=2 IA=32.0588  IB=66.8991
!Ic=98.4347  Ir=0.549  ROSYM=3  V(3)=~760. cm-1  Nu=3227,3209,3198,3185,3173,
!3168,3116,3055,3008,1633,1628,1504,1488,1476,1443,1438,1433,1387,1376,1312,1287,
!1211,1186,1168,1102,1081,1036,1033,1019,987,952.950,895,876,863,794,765,756,733,
!692,602,560,557,524,459,421,312,228,209,144  HF298=62.7 kcal  REF=Lifshitz
!Dubnikova JPC A 108,(2004),3430  DFT QCISD(T)//B3LYP/(cc-pVDZ) calc
!{HF298=60.264 kcal  REF=MOPAC 2000 PM3}  Max Lst Sq Error Cp @ 200 K 0.73%.
!C10H9 1-methyl    A03/05C 10.H  9.   0.   0.G   200.000  6000.000  B 129.17846 1
! 1.90083931E+01 3.18459404E-02-1.15126596E-05 1.86706540E-09-1.12145139E-13    2
! 2.23250010E+04-7.80332683E+01 4.07035729E-01 4.80530672E-02 6.13610491E-05    3
!-1.25042167E-07 5.63176095E-11 2.89729160E+04 2.60120139E+01 3.15516849E+04    4
!862559-83-9
!C10H9  2-Hydro-Naphthalene Radical   STATWT = 2   Ia = 27.990458  Ib = 71.911452
!Ic = 99.39347  NU= 3126,3110,3106,3095,3093,3090,3082,2851,2843,1636,1575,1528,
!1473,1430,1416,1397,1375,1353,1319,1260,1218,1185,1150,1137,1135,1112,1029,1016,
!949,928,900,899,891,886,831,764,761,734(2),678,667,594,525,491,484,445,390,344,
!256,169,125.  REF =Curran et al, JPCRD 29,(2000),463    Hf(298)= 54.86 kcal/mole
!REF = Marinov et al, Comb. Sci. Technol. 116-117,(1996), 211.   Max Lst Sq Error
!Cp @ 200 K  0.87%
naphthyl2H    Rad T 7/98C 10.H  9.   0.   0.G   200.000  6000.000 3000.0       1
 1.96879334E+01 3.20520257E-02-1.16715110E-05 1.90182471E-09-1.14603906E-13    2
 1.80099777E+04-8.29833882E+01-1.21356342E+00 5.48913745E-02 5.55281159E-05    3
-1.24860759E-07 5.75105005E-11 2.52575495E+04 3.28077928E+01 2.76064663E+04    4
! copy from C10H8
C6H4C2HC2H3             C  10H   8          G    300.00   4000.00 1401.00      1
 .234023214E+02 .242434427E-01-.836282016E-05 .130620111E-08-.761153748E-13    2
 .651941329E+04-.107433208E+03-.883645988E+01 .109300567E+00-.955200914E-04    3
 .421647669E-07-.739851710E-11 .166533366E+05 .621064766E+02                   4
!benzofulvenyl c10h7  assume naphthyl
Benzofulvenyl           C  10H   7          G    300.00   4000.00 1000.00      1
 .146529084E+02 .356159360E-01-.121796480E-04 .138747960E-08 .000000000E+00    2
 .405898415E+05-.575649187E+02-.631700500E+01 .913910790E-01-.608201990E-04    3
 .152228010E-07 .000000000E+00 .464268700E+05 .512234700E+02                   4
! copy from C10H8
C6H5CHCHCCH             C  10H   8          G    300.00   4000.00 1401.00      1
 .234023214E+02 .242434427E-01-.836282016E-05 .130620111E-08-.761153748E-13    2
 .651941329E+04-.107433208E+03-.883645988E+01 .109300567E+00-.955200914E-04    3
 .421647669E-07-.739851710E-11 .166533366E+05 .621064766E+02                   4
! to connect
C6H4CH3        RadT10/13C  7.H  7.   0.   0.G   200.000  6000.000 3000.00      1
 1.28543060E+01 2.42712778E-02-8.75277064E-06 1.41703290E-09-8.50082345E-14    2
 3.10872386E+04-4.29177096E+01 2.43474215E+00 2.10368651E-02 7.20305506E-05    3
-1.14038924E-07 4.82416036E-11 3.53949018E+04 1.83045052E+01 3.74896416E+04    4
C7H6         G3SX B3LYPTC   7H   6    0    0G   300.000  5000.000 1401.00      1
 1.70564548E+01 1.67766601E-02-5.75637904E-06 8.95748927E-10-5.20574674E-14    2
 3.43929834E+04-6.83510071E+01-3.96406850E+00 7.40750426E-02-6.68009279E-05    3
 3.06821623E-08-5.59258820E-12 4.08575050E+04 4.16088550E+01                   4
C7H5         G3SX ref819C   7H   5    0    0G   300.000  5000.000 1404.00      1
 1.65644050E+01 1.44569152E-02-4.91369020E-06 7.59739947E-10-4.39556749E-14    2
 4.96364603E+04-6.29487260E+01-2.77567748E+00 6.97210344E-02-6.63891369E-05    3
 3.18329494E-08-5.98040634E-12 5.53261073E+04 3.73111448E+01                   4  
CYC5H4                  C   5H   4          G    200.00   3500.00 1310.00      1
 6.52292919e+00 1.75112106e-02-7.24525264e-06 1.36814029e-09-9.77801928e-14    2
 6.01459587e+04-1.09295466e+01-1.67820638e+00 4.25528459e-02-3.59188809e-05    3
 1.59603175e-08-2.88254684e-12 6.22946562e+04 3.08507210e+01                   4
C5H3               20387C   5H   3          G  0300.00   5000.00  1000.00      1
 0.01078762E+03 0.09539619E-01-0.03206745E-04 0.04733323E-08-0.02512135E-12    2
 0.06392904E+06-0.03005444E+03 0.04328720E+02 0.02352480E+00-0.05856723E-04    3
-0.01215449E-06 0.07726478E-10 0.06588531E+06 0.04173259E+02                   4
C5H2               20587C   5H   2          G  0300.00   5000.00  1000.00      1
 0.01132917E+03 0.07424057E-01-0.02628189E-04 0.04082541E-08-0.02301333E-12    2
 0.07878706E+06-0.03617117E+03 0.03062322E+02 0.02709998E+00-0.01009170E-03    3
-0.01272745E-06 0.09167219E-10 0.08114969E+06 0.07071078E+02                   4
C5H5CH3                 C   6H   8          G    300.00   5000.00 1399.00      1
 .154352848E+02 .199801707E-01-.680270423E-05 .105349633E-08-.610336727E-13    2 
 .447456576E+04-.636393642E+02-.665320026E+01 .744640477E-01-.582864186E-04    3 
 .231603543E-07-.369017129E-11 .117669311E+05 .538162769E+02                   4
C7H7O2     QB3-MF11    0C   7H   7O   2    0G   300.00   5000.00  1000.00      1   
 1.71115179E+01 2.68198282E-02-1.06205723E-05 1.91920856E-09-1.30061244E-13    2
 6.71623207E+03-6.12436900E+01-2.24622429E+00 7.26022303E-02-3.67327921E-05    3
-8.74034681E-09 1.01564683E-11 1.24729027E+04 4.07042530E+01                   4
O2C6H4CH3    9/21/15    C   7H   7O   2    0G   300.000  5000.000 1408.000    21
 2.12862164E+01 1.93020680E-02-6.48485440E-06 9.95146950E-10-5.72828260E-14    2
 3.19865442E+03-8.60791351E+01-5.17635366E+00 9.32722534E-02-8.64517889E-05    3
 4.02042133E-08-7.33445923E-12 1.10698763E+04 5.15568699E+01                   4
OC6H4CH2          012508C   7H   6O   1     G   300.000  5000.000 1000.00      1
 1.24204756E+01 2.70171830E-02-1.09476851E-05 2.02705529E-09-1.40757462E-13    2
 4.49159466E+02-4.10236260E+01-6.21979546E-01 5.14918065E-02-6.11682462E-06    3
-2.88887155E-08 1.45119845E-11 4.44241036E+03 2.88224802E+01                   4
C6H5CH2O   4/14/94 THE.MC   7H   7O   1    0G   300.000  5000.000 1392.000     1
 1.78843033E+01 2.09011735E-02-7.21832713E-06 1.12839851E-09-6.57955260E-14    2
 4.93182818E+03-7.01304667E+01-4.77736690E+00 7.51049308E-02-5.68532831E-05    3
 2.18290029E-08-3.38134298E-12 1.26234438E+04 5.10429366E+01                   4
BZCOOH                  C   7H   8O   2    0G   300.000  5000.000 1388.000    31
 2.32849942E+01 2.11249905E-02-7.42176803E-06 1.17341778E-09-6.89572814E-14    2
-1.39352842E+04-9.56328725E+01-3.90619768E+00 8.82323518E-02-7.17190897E-05    3
 2.95644635E-08-4.91898930E-12-4.87198921E+03 4.90970451E+01                   4
C6H5O2                  H  5 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! LPM DHof 32.27 from automech C6H5+O2 paper
 9.44965310E+00 3.18801989E-02-1.65680518E-05 4.14518064E-09-4.05117628E-13    2
 1.22263498E+04-2.37678892E+01 1.27515227E+00 3.32184432E-02 4.35123037E-05    3
-9.12211721E-08 4.17171362E-11 1.51220807E+04 2.25793608E+01                   4
C5H4OCHO                H  5 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! LPM DHof -10.59 from automech C6H5+O2 paper
 1.00985212E+01 3.12036079E-02-1.62342321E-05 4.06249384E-09-3.96944018E-13    2
-1.21349626E+04-2.43033607E+01 2.38805714E+00 3.67187218E-02 2.50017851E-05    3
-6.72167921E-08 3.18416750E-11-9.55529680E+03 1.85256231E+01                   4
OXEPINOXY               H  5 C  6 O  2 N  0 G    200.0    3000.0   1000.0      1    ! LPM DHof -10.46 from automech C6H5+O2 paper
 8.86498881E+00 3.32321836E-02-1.72906475E-05 4.32839584E-09-4.23118854E-13    2
-1.20117732E+04-1.97833766E+01 1.10410411E+00 3.78525311E-02 2.71779716E-05    3
-7.06186149E-08 3.31958100E-11-9.37096841E+03 2.35498633E+01                   4
C6H5CO                  C   7H   5O   1    0G   300.000  5000.000 1396.000    11
 1.79587471E+01 1.58218495E-02-5.48154854E-06 8.58709339E-10-5.01435299E-14    2
 3.78486787E+03-7.06341032E+01-1.71526142E+00 6.53320500E-02-5.36914036E-05    3
 2.23697440E-08-3.73946626E-12 1.02136508E+04 3.36880709E+01                   4
RBBENZOOH  3/19/ 9 THERMC  14H  14O   2    0G   300.000  5000.000 1395.000    51
 4.01427062E+01 3.93395367E-02-1.37664348E-05 2.17056135E-09-1.27304368E-13    2
-1.39277882E+04-1.84904308E+02-1.04261530E+01 1.68709899E-01-1.42892982E-04    3
 6.15601039E-08-1.06485940E-11 2.47291567E+03 8.26365480E+01                   4
RBBENZOO   3/19/ 9 THERMC  14H  13O   2    0G   300.000  5000.000 1394.000    41
 3.76701265E+01 3.91886728E-02-1.36838688E-05 2.15430957E-09-1.26216113E-13    2
 4.38748283E+03-1.69872607E+02-9.53800906E+00 1.60095043E-01-1.34982895E-04    3
 5.84090458E-08-1.01919995E-11 1.97390228E+04 7.99308597E+01                   4
QBBENZOOH  3/19/ 9 THERMC  14H  13O   2    0G   300.000  5000.000 1394.000    41
 4.02968908E+01 3.71210431E-02-1.30088643E-05 2.05309245E-09-1.20495552E-13    2
 3.67900543E+03-1.86479334E+02-8.32529422E+00 1.61762848E-01-1.37724101E-04    3
 5.95672829E-08-1.03363053E-11 1.94259748E+04 7.06782085E+01                   4
ZBBENZ        9/ 9 THERMC  14H  13O   4    0G   300.000  5000.000 1391.000    71
 4.48785960E+01 3.75685709E-02-1.32824040E-05 2.10858085E-09-1.24255944E-13    2
-9.97231472E+03-2.04041648E+02-9.40646930E+00 1.77878119E-01-1.55260847E-04    3
 6.84418245E-08-1.20655066E-11 7.52457116E+03 8.27128410E+01                   4
KHYBBENZ     19/ 9 THERMC  14H  12O   3    0G   300.000  5000.000 1393.000    41
 4.03057402E+01 3.72594407E-02-1.30902950E-05 2.06942373E-09-1.21596482E-13    2
-2.78034193E+04-1.82398868E+02-7.77794671E+00 1.57347464E-01-1.29564931E-04    3
 5.40605490E-08-9.07699935E-12-1.19364337E+04 7.29984559E+01                   4
C14H13O    3/19/ 9 THERMC  14H  13O   1    0G   300.000  5000.000 1397.000    31
 3.62205336E+01 3.75634484E-02-1.29678295E-05 2.02688785E-09-1.18180078E-13    2
 5.74597621E+03-1.65590808E+02-1.19190739E+01 1.59861239E-01-1.33105430E-04    3
 5.60228564E-08-9.42896323E-12 2.13328544E+04 8.92151705E+01                   4
BZCOOH                  C   7H   8O   2    0G   300.000  5000.000 1388.000    31
 2.32849942E+01 2.11249905E-02-7.42176803E-06 1.17341778E-09-6.89572814E-14    2
-1.39352842E+04-9.56328725E+01-3.90619768E+00 8.82323518E-02-7.17190897E-05    3
 2.95644635E-08-4.91898930E-12-4.87198921E+03 4.90970451E+01                   4
RBBENZ                  C  14H  13          G    300.00   4000.00 1000.00      1
 .299291000E+02 .383042200E-01-.118663300E-04 .177305900E-08-.104476700E-12    2
 .197099600E+05-.131713300E+03-.766215500E+01 .133505200E+00-.973103200E-04    3
 .342829900E-07-.478937100E-11 .309915700E+05 .658134800E+02                   4
STILB                   C  14H  12          G    300.00   4000.00 1000.00      1
 .268497500E+02 .428429300E-01-.150785000E-04 .246643600E-08-.154717900E-12    2
 .164217700E+05-.117418300E+03-.792701200E+01 .132075300E+00-.881173300E-04    3
 .190952300E-07 .176879600E-11 .263867200E+05 .640743300E+02                   4
C14H12O   10/19/15      C  14H  12O   1    0G   300.000  5000.000 1394.000    31 
 3.48141204E+01 3.67953648E-02-1.28282619E-05 2.01783856E-09-1.18158524E-13    2
-1.68668837E+04-1.61938007E+02-9.56374055E+00 1.44801295E-01-1.13794706E-04    3
 4.50882665E-08-7.17648586E-12-2.00559523E+03 7.46678724E+01                   4
!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
!************************BUTANOIC ACID SET **************************************!
!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
C3H7COOH   ButAcidT12/07C  4.H  8.O  2.   0.G   200.000  6000.000 1000.        1   !Burcat
 1.04116580E+01 2.47964316E-02-8.90592565E-06 1.43428158E-09-8.56419203E-14    2
-6.01225120E+04-2.47412226E+01 6.55568876E+00 1.19881222E-03 9.25041110E-05    3
-1.19593964E-07 4.69861556E-11-5.74283767E+04 3.36226959E+00-5.48174043E+04    4
CH2COOH                 C   2H   3O   2     G  0300.000  5000.000 1000.        1 !Thergas
 0.93029661E+01 0.69815558E-02-0.17180930E-05 0.21747887E-09-0.11452205E-13    2
-0.33653477E+05-0.23130653E+02 0.12598374E+00 0.34687348E-01-0.34489818E-04    3
 0.18876753E-07-0.44256933E-11-0.31187451E+05 0.23825567E+02                   4
CH2CH2COOH              C   3H   5O   2     G  0300.00   5000.00  1000.00      1 !Thergas
 0.13256764E+02 0.88558299E-02-0.20110283E-05 0.23953006E-09-0.12087953E-13    2
-0.34287797E+05-0.40638344E+02-0.21509118E+01 0.64166412E-01-0.84363666E-04    3
 0.58959127E-07-0.16281953E-10-0.30510459E+05 0.36154118E+02                   4
RBUTANOICB              C   4H   7O   2     G  0300.00   5000.00  1000.00      1        !sec beta pentanoic, needed better estimate
 0.17189188E+02 0.20083707E-01-0.55279124E-05 0.75932416E-09-0.42271813E-13    2
-0.42307125E+05-0.57420525E+02-0.27705753E+01 0.90017982E-01-0.10568813E-03    3
 0.69284084E-07-0.18381326E-10-0.37391141E+05 0.42345650E+02                   4
RBUTANOICA              C   4H   7O   2     G  0300.00   5000.00  1000.00      1        !sec alfa pentanoic, needed better estimate
 0.17195915E+02 0.21016909E-01-0.60015391E-05 0.84707413E-09-0.48064749E-13    2
-0.44621500E+05-0.60233444E+02-0.23888919E+01 0.86213857E-01-0.93720431E-04    3
 0.57221794E-07-0.14316034E-10-0.39635621E+05 0.38491531E+02                   4
RBUTANOICC              C   4H   7O   2     G  0300.00   5000.00  1000.00      1        !prim  pentanoic, needed better estimate
 0.17552582E+02 0.20030502E-01-0.55556238E-05 0.76777634E-09-0.42941223E-13    2
-0.41376172E+05-0.59720062E+02-0.25150366E+01 0.87286346E-01-0.96496748E-04    3
 0.59345126E-07-0.14867392E-10-0.36302215E+05 0.41297184E+02                   4
C2H5CHCO                C   4H   6O   1    0G   200.000  6000.000 1000.000    21    !from Burcat
 1.12344400E+01 1.66857869E-02-5.99141532E-06 9.66147739E-10-5.78333791E-14    2
-1.89013763E+04-3.34159921E+01 2.98852451E+00 2.04971182E-02 3.56246580E-05    3
-6.38395109E-08 2.75663362E-11-1.57565701E+04 1.36212503E+01-1.37529115E+04    4
C3H7CHCO                C   5H   8O   1    0G   200.000  6000.000 1000.000    21    !corrected group additivity burcat
 1.50903576E+01	1.96657858E-02-6.48018243E-06 9.27416519E-10-4.70728721E-14    2
-2.31212013E+04-5.24144550E+01 3.54009480E-01 5.33779762E-02-2.80581975E-05    3
 2.90860000E-12	3.47960790E-12-1.85224858E+04 2.58839478E+01                   4
C3H5COOH-1              C   4H   6O   2     G  0200.00   6000.00  1000.00      1   !Burcat
 1.25067898E+01 1.79507069E-02-6.45643374E-06 1.04141105E-09-6.22628191E-14    2
-4.92096261E+04-3.74168332E+01 3.40323244E+00 2.69846381E-02 2.63698041E-05    3
-5.87466892E-08 2.69692257E-11-4.60243863E+04 1.31927575E+01-4.36807162E+04    4
C2H3COOH                C   3H   4O   2     G  0200.00   6000.00  1000.00      1   !Burcat
 1.04962923E+01 1.20559957E-02-4.34149310E-06 6.99425892E-10-4.18003976E-14    2
-4.37332461E+04-2.75425657E+01 1.24227207E+00 3.00698605E-02-1.48206586E-06    3
-2.42738150E-08 1.33121686E-11-4.08667843E+04 2.19242842E+01-3.92146683E+04    4
CH2COOH                 C   2H   3O   2     G  0300.00   5000.00  1000.00      1
 0.93029661E+01 0.69815558E-02-0.17180930E-05 0.21747887E-09-0.11452205E-13    2
-0.33653477E+05-0.23130653E+02 0.12598374E+00 0.34687348E-01-0.34489818E-04    3
 0.18876753E-07-0.44256933E-11-0.31187451E+05 0.23825567E+02                   4
CH2CH2COOH              C   3H   5O   2     G  0300.00   5000.00  1000.00      1
-0.63459964E+01 0.40684473E-01-0.16808332E-04 0.30763088E-08-0.20875162E-12    2
-0.26339281E+05 0.69442528E+02-0.12847569E+01 0.57524763E-01-0.66488785E-04    3
 0.38840408E-07-0.82382261E-11-0.30595645E+05 0.32566666E+02                   4
!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
!************************PENTANOIC ACID SET *************************************!
!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
C4H9COOH                C   5H  10O   2     G  0300.00   5000.00  1000.00      1
 0.13259649E+02 0.30104950E-01-0.10327794E-04 0.16574947E-08-0.10252313E-12    2
-0.64599336E+05-0.38116192E+02-0.14140378E+01 0.76504208E-01-0.63748710E-04    3
 0.27372781E-07-0.41224650E-11-0.60943137E+05 0.35990471E+02                   4
RPENTANOICB             C   5H   9O   2     G  0300.00   5000.00  1000.00      1        !sec beta pentanoic THERGAS
 0.17189188E+02 0.20083707E-01-0.55279124E-05 0.75932416E-09-0.42271813E-13    2
-0.42307125E+05-0.57420525E+02-0.27705753E+01 0.90017982E-01-0.10568813E-03    3
 0.69284084E-07-0.18381326E-10-0.37391141E+05 0.42345650E+02                   4
RPENTANOICA             C   5H   9O   2     G  0300.00   5000.00  1000.00      1        !sec alfa pentanoic THERGAS
 0.17195915E+02 0.21016909E-01-0.60015391E-05 0.84707413E-09-0.48064749E-13    2
-0.44621500E+05-0.60233444E+02-0.23888919E+01 0.86213857E-01-0.93720431E-04    3
 0.57221794E-07-0.14316034E-10-0.39635621E+05 0.38491531E+02                   4
RPENTANOICC             C   5H   9O   2     G  0300.00   5000.00  1000.00      1        !sec gam
 0.16945580E+02 0.20560963E-01-0.57434822E-05 0.79954027E-09-0.45031782E-13    2
-0.42261293E+05-0.56176674E+02-0.16730661E+01 0.82255505E-01-0.88211753E-04    3
 0.53189538E-07-0.13042655E-10-0.37498469E+05 0.37762043E+02                   4
RPENTANOICD             C   5H   9O   2     G  0300.00   5000.00  1000.00      1        !prim  pentanoic, THERGAS
 0.17552582E+02 0.20030502E-01-0.55556238E-05 0.76777634E-09-0.42941223E-13    2
-0.41376172E+05-0.59720062E+02-0.25150366E+01 0.87286346E-01-0.96496748E-04    3
 0.59345126E-07-0.14867392E-10-0.36302215E+05 0.41297184E+02                   4
C4H7COOH-1              C   5H   8O   2     G  0300.00   5000.00  1000.00      1
 1.45172873E+01	2.38454181E-02-8.57137438E-06 1.38339621E-09-8.27252406E-14    2
-5.46860061E+04-4.72911007E+01 5.56419281E+00 2.38994157E-02 5.42216741E-05    3
-9.32195634E-08	4.06262828E-11-5.11819883E+04 4.46123080E+00                   4
!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
!!!!!!!!!!!!!!! Heufer et al. Lumped nC3-C6 alcohols cyclic ethers!!!!!!!!!!!!!!!!
C6OHCYETH    11    THERMC   6H  12O   2    0G   300.000  5000.000 1397.000    11
 1.87792328E+01 2.52510031E-02-8.71951941E-06 1.36261690E-09-7.94233655E-14    2
-5.98486874E+04-8.02952910E+01-5.28245732E+00 8.05420193E-02-5.65771489E-05    3
 1.99013096E-08-2.79015119E-12-5.14625083E+04 4.91527811E+01                   4
C5OHCYETH    11    THERMC   5H  10O   2    0G   300.000  5000.000 1397.000    11
 1.87792328E+01 2.52510031E-02-8.71951941E-06 1.36261690E-09-7.94233655E-14    2
-5.98486874E+04-8.02952910E+01-5.28245732E+00 8.05420193E-02-5.65771489E-05    3
 1.99013096E-08-2.79015119E-12-5.14625083E+04 4.91527811E+01                   4
C4OHCYETH   5/6/11 THERMC   4H   8O   2    0G   300.000  5000.000 1401.000    21
 1.53974801E+01 1.99867721E-02-6.88756825E-06 1.07490272E-09-6.25966766E-14    2
-5.33539148E+04-5.82489337E+01-4.33894975E+00 6.58008223E-02-4.69211010E-05    3
 1.67037853E-08-2.35942205E-12-4.65427473E+04 4.77300998E+01                   4
C3OHCYETH   5/6/11 THERMC   3H   6O   2    0G   200.000  6000.000 1000.000    21
 1.03094493E+01 1.72095929E-02-6.11612099E-06 9.80636991E-10-5.84379268E-14    2
-3.36703047E+04-2.78187504E+01 3.21008917E+00 1.25973594E-02 5.89962103E-05    3
-9.09895491E-08 3.85110105E-11-3.06902814E+04 1.42923264E+01-2.88136831E+04    4	
!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
!*******************************************************************************!
!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
!NOx MODULE (from Burcat http://garfield.chem.elte.hu/Burcat/THERM.DAT)
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NO                RUS 89N   1O   1    0    0G   200.000  6000.000 1000.        1
 3.26071234E+00 1.19101135E-03-4.29122646E-07 6.94481463E-11-4.03295681E-15    2
 9.92143132E+03 6.36900518E+00 4.21859896E+00-4.63988124E-03 1.10443049E-05    3
-9.34055507E-09 2.80554874E-12 9.84509964E+03 2.28061001E+00 1.09770882E+04    4
N2O               L 7/88N   2O   1    0    0G   200.000  6000.000 1000.        1
 0.48230729E+01 0.26270251E-02-0.95850872E-06 0.16000712E-09-0.97752302E-14    2
 0.80734047E+04-0.22017208E+01 0.22571502E+01 0.11304728E-01-0.13671319E-04    3
 0.96819803E-08-0.29307182E-11 0.87417746E+04 0.10757992E+02 0.98141682E+04    4
NO2               L 7/88N   1O   2    0    0G   200.000  6000.000 1000.        1
 0.48847540E+01 0.21723955E-02-0.82806909E-06 0.15747510E-09-0.10510895E-13    2
 0.23164982E+04-0.11741695E+00 0.39440312E+01-0.15854290E-02 0.16657812E-04    3
-0.20475426E-07 0.78350564E-11 0.28966180E+04 0.63119919E+01 0.41124701E+04    4
HNO               ATcT/AH  1.N  1.O  1.   0.G   200.000  6000.000 1000.        1
 3.16598124E+00 2.99958892E-03-3.94376786E-07-3.85344089E-11 7.07602668E-15    2
 1.17726311E+04 7.64511172E+00 4.53525574E+00-5.68543377E-03 1.85198540E-05    3
-1.71881225E-08 5.55818157E-12 1.16183003E+04 1.74315886E+00 1.28500657E+04    4
HNNO                    H   1O   1N   2     G    300.00   4000.00 1500.00      1 ! Not present in Burcat. Old Thermochemistry data were kept
 .699121930E+01 .187597000E-02-.212458400E-06-.671047200E-10 .123050800E-13    2
 .249756641E+05-.112352384E+02 .223829800E+01 .135920000E-01-.117987300E-04    3
 .539297100E-08-.101085900E-11 .266025900E+05 .141367900E+02                   4
!HNO2 equil  ATcT  T 9/11H  1.N  1.O  2.   0.G   200.000  6000.000 1000.        1
! 5.79182717E+00 3.65162554E-03-1.29293390E-06 2.06892796E-10-1.23154749E-14    2
!-1.15953895E+04-4.05538852E+00 3.21415915E+00 8.12778066E-03 1.65998916E-06    3
!-9.52814708E-09 4.87131424E-12-1.07830727E+04 9.82200056E+00-9.46538040E+03    4
HNO2              ATcT3EH   1N   1O   2    0G    200.00   6000.00 1000.00      1 ! Glarborg PECS 2018
 4.66358504E+00 4.89854351E-03-1.79694193E-06 2.94420361E-10-1.78235577E-14    2
-7.25216334E+03-3.06053640E-02 4.03779347E+00-4.46123109E-03 3.19440815E-05    3
-3.79359490E-08 1.44570885E-11-6.53088236E+03 5.90620097E+00-5.31122753E+03    4
HONO              ATcT3EH   1N   1O   2    0G    200.00   6000.00 1000.00      1 ! Glarborg PECS 2018
 5.79144641E+00 3.64630732E-03-1.29112765E-06 2.06498233E-10-1.22138679E-14    2
-1.15974343E+04-4.07145349E+00 3.16416438E+00 8.50517773E-03 5.48561573E-07    3
-8.27656474E-09 4.39957151E-12-1.07744086E+04 1.00231941E+01-9.46242812E+03    4
HONO2             T 8/03H  1.N  1.O  3.   0.G   200.000  6000.000 1000.        1 ! Is HNO3 in Burcat database
 8.03098942E+00 4.46958589E-03-1.72459491E-06 2.91556153E-10-1.80102702E-14    2
-1.93138183E+04-1.62616537E+01 1.69329154E+00 1.90167702E-02-8.25176697E-06    3
-6.06113827E-09 4.65236978E-12-1.74198909E+04 1.71839838E+01-1.61524852E+04    4
N2H2 equil & transT 9/11N  2.H  2.   0.   0.G   200.000  6000.000 1000.        1
 1.31115117E+00 9.00187208E-03-3.14911824E-06 4.81449581E-10-2.71897891E-14    2
 2.33863341E+04 1.64091067E+01 4.91066031E+00-1.07791880E-02 3.86516489E-05    3
-3.86501698E-08 1.34852134E-11 2.28241901E+04 9.10273396E-02 2.40806734E+04    4
H2NN Isodiazene   T 9/11N  2.H  2.   0.   0.G   200.000  6000.000 1000.        1 ! Is 'N2H2 Isodiazene' in Burcat database
 3.05903670E+00 6.18382347E-03-2.22171165E-06 3.58539206E-10-2.14532905E-14    2
 3.48530149E+04 6.69893515E+00 4.53204001E+00-7.32418578E-03 3.00803713E-05    3
-3.04000551E-08 1.04700639E-11 3.49580003E+04 1.51074195E+00 3.61943157E+04    4
HNNO      5/30/18 THERM N  2.H  1.O  1    0.G   300.000  5000.000 1790.000    61 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 2.15594002E+06-4.13111192E+03 2.65627771E+00-6.70395293E-04 5.57827338E-08    2
-8.03468100E+08-1.18702032E+07-8.96779017E-01 3.69714359E-02-4.80099825E-05    3
 2.62274393E-08-5.11382966E-12 2.68675048E+04 2.64521806E+01                   4
NH2NO     5/30/18 THERM N  2.H  2.O  1    0.G   300.000  5000.000 1371.000    61 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 7.93898100E+00 5.21842622E-03-2.12493130E-06 3.53331059E-10-2.12447889E-14    2
 5.42322972E+03-1.84299492E+01 1.85914077E+00 1.68525394E-02-9.37240888E-06    3
 1.71380329E-09 4.84625807E-14 7.78108234E+03 1.51172833E+01                   4
HNOH trans & Equ  T11/11H  2.N  1.O  1.   0.G   200.000  6000.000 1000.        1
 3.98321933E+00 4.88846374E-03-1.65086637E-06 2.55371446E-10-1.48308561E-14    2
 1.05780106E+04 3.62582838E+00 3.95608248E+00-3.02611020E-03 2.56874396E-05    3
-3.15645120E-08 1.24084574E-11 1.09199790E+04 5.55950983E+00 1.21354115E+04    4
NH2OH             ATcT/AN  1.H  3.O  1.   0.G   200.000  6000.000 1000.        1
 3.88112502E+00 8.15708448E-03-2.82615576E-06 4.37930933E-10-2.52724604E-14    2
-6.86018419E+03 3.79156136E+00 3.21016092E+00 6.19671676E-03 1.10594948E-05    3
-1.96668262E-08 8.82516590E-12-6.58148481E+03 7.93293571E+00-5.28593988E+03    4
NH3               ATcT3EH   3N   1    0    0G    200.00   4000.00 1000.00      1 ! Glarborg PECS 2018
 2.36074311E+00 6.31850146E-03-2.28966806E-06 4.11767411E-10-2.90836787E-14    2
-6.41596473E+03 8.02154329E+00 4.14027871E+00-3.58489142E-03 1.89475904E-05    3
-1.98833970E-08 7.15267961E-12-6.68545158E+03-1.66754883E-02-5.47888720E+03    4
N2H4 HYDRAZINE    L 5/90N   2H   4    0    0G   200.000  6000.000 1000.        1
 4.93957357E+00 8.75017187E-03-2.99399058E-06 4.67278418E-10-2.73068599E-14    2
 9.28265548E+03-2.69439772E+00 3.83472149E+00-6.49129555E-04 3.76848463E-05    3
-5.00709182E-08 2.03362064E-11 1.00893925E+04 5.75272030E+00 1.14474575E+04    4
HCN               ATcT/AH  1.C  1.N  1.   0.G   200.000  6000.000 1000.        1
 3.80231648E+00 3.14630087E-03-1.06315727E-06 1.66185438E-10-9.79891962E-15    2
 1.42849502E+04 1.57501632E+00 2.25901199E+00 1.00510475E-02-1.33514567E-05    3
 1.00920479E-08-3.00880408E-12 1.45903166E+04 8.91631960E+00 1.56111424E+04    4
HNC               ATcT/AH  1.N  1.C  1.   0.G   200.000  6000.000 1000.        1
 4.22248262E+00 2.59458082E-03-8.58480324E-07 1.30744940E-10-7.50339813E-15    2
 2.17156730E+04-7.79706410E-02 2.30186822E+00 1.54157449E-02-3.13261898E-05    3
 3.08816218E-08-1.11912204E-11 2.19306327E+04 8.14749128E+00 2.30810956E+04    4
HNCO Isocyanic AciA 5/05H  1.N  1.C  1.O  1.G   200.000  6000.000 1000.        1
 5.30045051E+00 4.02250821E-03-1.40962280E-06 2.23855342E-10-1.32499966E-14    2
-1.61995274E+04-3.11770684E+00 2.24009031E+00 1.45600497E-02-1.54352330E-05    3
 8.55535028E-09-1.79631611E-12-1.54589951E+04 1.21663775E+01-1.42642740E+04    4
HCNO Fulminic AcidA 5/05H  1.N  1.C  1.O  1.G   200.000  6000.000 1000.        1
 5.91979744E+00 4.00114600E-03-1.42063343E-06 2.27569621E-10-1.35504870E-14    2
 1.80385534E+04-8.26935223E+00 6.07949401E-01 2.82182431E-02-4.60451618E-05    3
 3.82559486E-08-1.23226501E-11 1.90714209E+04 1.69199098E+01 2.01698706E+04    4
HOCN Cyanic Acid  A 5/05H  1.N  1.C  1.O  1.G   200.000  6000.000 1000.        1
 5.28767714E+00 4.01746511E-03-1.40407465E-06 2.22562614E-10-1.31562375E-14    2
-3.77409807E+03-2.64470976E+00 2.88943546E+00 1.16487242E-02-1.08005006E-05    3
 5.44138776E-09-1.06857286E-12-3.15296691E+03 9.51295652E+00-1.85890558E+03    4
CH3NO NitrosomethyT12/09C  1.H  3.N  1.O  1.G   200.000  6000.000 1000.        1
 5.04711802E+00 9.21544305E-03-3.29034831E-06 5.28940397E-10-3.15689858E-14    2
 6.23718102E+03-7.74395570E-01 5.18534727E+00-6.34085575E-03 4.57171139E-05    3
-5.30421813E-08 1.99501601E-11 6.93771506E+03 2.18492659E+00 8.51040025E+03    4
CH3NO2            T01/00C   1H   3N   1O   2G   200.000  6000.000 1000.        1
 6.73034758E+00 1.09601272E-02-4.05357875E-06 6.67102246E-10-4.04686823E-14    2
-1.29143475E+04-1.01800883E+01 3.54053638E+00 1.86559899E-03 4.44946580E-05    3
-5.87057133E-08 2.30684496E-11-1.11385976E+04 1.06884657E+01-9.71208165E+03    4
CH3ONO            A 5/05C  1.H  3.O  2.N  1.G   200.000  6000.000 1000.        1
 6.93605239E+00 9.97319424E-03-3.60642537E-06 5.83462161E-10-3.50058729E-14    2
-1.08381899E+04-6.98144573E+00 6.15261387E+00-2.91937431E-03 4.14526828E-05    3
-4.93954776E-08 1.85608328E-11-9.85260262E+03 8.04057190E-01-7.87057806E+03    4
CH3ONO2           T05/98C   1H   3N   1O   3G   200.000  6000.000 1000.        1
 9.77845489E+00 1.10069541E-02-4.25928645E-06 7.18198185E-10-4.42041793E-14    2
-1.88804487E+04-2.39163197E+01 3.91363583E+00 1.52137945E-02 1.73479131E-05    3
-3.37074473E-08 1.44322204E-11-1.66103232E+04 9.44208392E+00-1.46737980E+04    4
CH3CN Methyl-Cya  T01/03C  2.H  3.N  1.   0.G   200.000  6000.000 1000.        1
 5.09921882E+00 9.69585649E-03-3.48051966E-06 5.61420173E-10-3.35835856E-14    2
 6.60967324E+03-3.36087178E+00 3.82392803E+00 4.08201943E-03 2.16209537E-05    3
-2.89807789E-08 1.12962700E-11 7.44430382E+03 5.52656156E+00 8.90492212E+03    4
N                 L 6/88N   1    0    0    0G   200.000  6000.000 1000.        1
 0.24159429E+01 0.17489065E-03-0.11902369E-06 0.30226244E-10-0.20360983E-14    2
 0.56133775E+05 0.46496095E+01 0.25000000E+01 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.56104638E+05 0.41939088E+01 0.56850013E+05    4
NO3               ATcT/AN  1.O  3.   0.   0.G   200.000  6000.000 1000.        1
 7.48347702E+00 2.57772064E-03-1.00945831E-06 1.72314063E-10-1.07154008E-14    2
 6.12990474E+03-1.41618136E+01 2.17359330E+00 1.04902685E-02 1.10472669E-05    3
-2.81561867E-08 1.36583960E-11 7.81290905E+03 1.46022090E+01 8.97563416E+03    4
NH                ATcT/AN  1.H  1.   0.   0.G   200.000  6000.000 1000.        1
 2.78372644E+00 1.32985888E-03-4.24785573E-07 7.83494442E-11-5.50451310E-15    2
 4.23461945E+04 5.74084863E+00 3.49295037E+00 3.11795720E-04-1.48906628E-06    3
 2.48167402E-09-1.03570916E-12 4.21059722E+04 1.84834973E+00 4.31525130E+04    4
NNH               T 8/11N  2.H  1.   0.   0.G   200.000  6000.000 1000.        1 ! Is N2H in Burcat database
 3.42744423E+00 3.23295234E-03-1.17296299E-06 1.90508356E-10-1.14491506E-14    2
 2.87676026E+04 6.39209233E+00 4.25474632E+00-3.45098298E-03 1.37788699E-05    3
-1.33263744E-08 4.41023397E-12 2.87932080E+04 3.28551762E+00 3.00058572E+04    4
NH2  AMIDOGEN RAD IU3/03N  1.H  2.   0.   0.G   200.000  3000.000 1000.        1
 2.59263049E+00 3.47683597E-03-1.08271624E-06 1.49342558E-10-5.75241187E-15    2
 2.15737320E+04 7.90565351E+00 4.19198016E+00-2.04602827E-03 6.67756134E-06    3
-5.24907235E-09 1.55589948E-12 2.11863286E+04-9.04785244E-02 2.23945849E+04    4
H2NO  RADICAL     T09/09N  1.H  2.O  1.   0.G   200.000  6000.000 1000.        1 ! From Glarborg thermo database (cannot find in Burcat)
 3.75555914E+00 5.16219354E-03-1.76387387E-06 2.75052692E-10-1.60643143E-14    2
 6.51826177E+03 4.30933053E+00 3.93201139E+00-1.64028165E-04 1.39161409E-05    3
-1.62747853E-08 6.00352834E-12 6.71178975E+03 4.58837038E+00 7.97044877E+03    4
N2H3   Rad.       T 7/11N  2.H  3.   0.   0.G   200.000  6000.000 1000.        1
 4.04483566E+00 7.31130186E-03-2.47625799E-06 3.83733021E-10-2.23107573E-14    2
 2.53241420E+04 2.88423392E+00 3.42125505E+00 1.34901590E-03 2.23459071E-05    3
-2.99727732E-08 1.20978970E-11 2.58198956E+04 7.83176309E+00 2.70438066E+04    4
CN                IU8/03C  1.N  1.   0.   0.G   200.000  6000.000 1000.        1
 3.39912850E+00 7.46548662E-04-1.41493852E-07 1.86747736E-11-1.26032540E-15    2
 5.16569715E+04 4.67148681E+00 3.61256069E+00-9.53015737E-04 2.13757271E-06    3
-3.05001808E-10-4.70518097E-13 5.17084034E+04 3.98238722E+00 5.27611901E+04    4
NCN  MethaneTetr  T 5/14C  1.N  2.   0.   0.G   200.000  6000.000 1000.        1
 5.68744173E+00 1.82662756E-03-7.07546249E-07 1.19515592E-10-7.31827071E-15    2
 5.15901177E+04-6.31954433E+00 2.79807977E+00 1.00008683E-02-9.59229469E-06    3
 4.75546842E-09-1.04340146E-12 5.24021705E+04 8.62129767E+00 5.36050832E+04    4
NCO  (NCO)        A 5/05N  1.C  1.O  1.   0.G   200.000  6000.000 1000.        1 ! Is CNO (NCO) in Burcat database
 5.08064474E+00 2.37443587E-03-9.07098904E-07 1.52286713E-10-9.31009234E-15    2
 1.35781204E+04-2.15734434E+00 2.77405177E+00 9.24523481E-03-9.91773586E-06    3
 6.68461303E-09-2.09520542E-12 1.42369570E+04 9.75458670E+00 1.53995606E+04    4
HNCN Cyanamide    T03/10C  1.H  1.N  2.   0.G   200.000  6000.000 1000.        1
 5.53846448E+00 3.89054126E-03-1.38104752E-06 2.21294765E-10-1.31827325E-14    2
 3.59635337E+04-3.39587098E+00 3.06754311E+00 1.06789939E-02-7.96224305E-06    3
 2.59883390E-09-1.27057612E-13 3.66623508E+04 9.41074995E+00 3.79863165E+04    4
H2CN  H2C=N*      T 1/11C  1.H  2.N  1.   0.G   200.000  6000.000 1000.        1 ! Is CH2N in Burcat database
 3.80315578E+00 5.47197362E-03-1.95314875E-06 3.13362403E-10-1.86249384E-14    2
 2.71302747E+04 3.31759436E+00 3.97799555E+00-3.43275801E-03 2.59134260E-05    3
-3.04692171E-08 1.16272717E-11 2.74854081E+04 4.43067396E+00 2.86930920E+04    4
C2N2 Dicyanogen   ATcT/AC  2.N  2.   0.   0.G   200.000  6000.000 1000.        1
 6.70549520E+00 3.64271185E-03-1.30939702E-06 2.16421413E-10-1.31193815E-14    2
 3.48824335E+04-1.04803146E+01 2.32928126E+00 2.61540993E-02-4.90009889E-05    3
 4.61923035E-08-1.64325831E-11 3.56900732E+04 9.86348075E+00 3.71976220E+04    4
CH2CN     1/16/17  THERMC  2.H  2.N  1.   0.G   300.000  5000.000 1414.000    61 ! K Sendt E Ikeda GB Bacskay JC Mackie JPCA 103 (1999) 1054-1072
 6.36314975E+00 6.36391885E-03-2.75175653E-06 5.78264246E-10-4.21050412E-14    2
 2.90725105E+04-8.80921516E+00 3.13213813E+00 1.42275608E-02-1.03390720E-05    3
 4.00717364E-09-6.45501720E-13 3.01853547E+04 8.46664206E+00                   4
HCNH  H*C=NH TransT11/11C  1.H  2.N  1.   0.G   200.000  6000.000 1000.        1
 4.04014700E+00 5.16591694E-03-1.82276828E-06 2.90299053E-10-1.71614589E-14    2
 3.11540211E+04 2.58894095E+00 3.97114555E+00-3.88875724E-03 2.92918950E-05    3
-3.57482411E-08 1.40303911E-11 3.15789298E+04 5.06388721E+00 3.27848544E+04    4
C3HN Cyano-Acety  A 2/05C  3.H  1.N  1.   0.G   200.000  6000.000 1000.        1
 7.44515032E+00 5.27107604E-03-1.86735278E-06 2.98683734E-10-1.77665376E-14    2
 4.16450237E+04-1.46187448E+01 5.87779106E-01 3.84323486E-02-6.61566501E-05    3
 5.72555769E-08-1.89892637E-11 4.29066005E+04 1.74909167E+01 4.43097371E+04    4
CH3NH2            T04/14C  1.H  5.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database (CH5N)
 4.46959661E+00 1.21969427E-02-4.31573211E-06 6.89638406E-10-4.09907834E-14    2
-4.86166208E+03-1.73983318E+00 4.93595327E+00-1.06687240E-02 6.66595644E-05    3
-7.68165338E-08 2.88891949E-11-3.96311166E+03 1.01955189E+00-2.51488061E+03    4
CH2NH             T 8/11C  1.H  3.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database (CH3N)
 3.44258358E+00 8.37600036E-03-2.97819078E-06 4.77352867E-10-2.84295062E-14    2
 8.97134621E+03 3.95595397E+00 4.79302577E+00-1.26841692E-02 5.69766521E-05    3
-6.34985251E-08 2.37023330E-11 9.41385818E+03 1.10277996E+00 1.06682174E+04    4
CH2NH2            T 8/11C  1.H  4.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database (*CH2NH2)
 4.55329728E+00 9.42002581E-03-3.20781399E-06 4.98961894E-10-2.90872284E-14    2
 1.58717284E+04-2.45945234E-02 2.85538164E+00 7.27364238E-03 1.65712636E-05    3
-2.70976978E-08 1.16327939E-11 1.66165986E+04 1.02444521E+01 1.78895690E+04    4
CH3NH             T03/10C  1.H  4.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database (CH3NH radical)
 4.02244380E+00 1.03512061E-02-3.64560169E-06 5.80491587E-10-3.44103829E-14    2
 1.95050854E+04 1.64483768E+00 4.70973738E+00-7.31946952E-03 4.95105509E-05    3
-5.72790480E-08 2.16523586E-11 2.00619432E+04 1.85460205E+00 2.14752744E+04    4
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
!PYRROLE MODULE
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
C4H5N     1/16/17  THERMC  4.H  5.N  1.   0.G   300.000  5000.000 1430.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 1.08130186E+01 1.48492978E-02-4.63893065E-06 6.75632087E-10-3.74350506E-14    2
 7.86128350E+03-3.62440836E+01-5.22833031E+00 6.28815185E-02-5.92617976E-05    3
 2.83624834E-08-5.27666016E-12 1.22545900E+04 4.59560293E+01                   4
C4H4N  Pyrridyl R T 7/14C  4.H  4.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database
 9.56455967E+00 1.37100337E-02-4.92563602E-06 7.95650357E-10-4.76637329E-14    2
 3.05922716E+04-2.78072307E+01 7.12951232E-01 1.73878483E-02 4.69371029E-05    3
-8.26955853E-08 3.67546269E-11 3.38297439E+04 2.23581694E+01 3.50837627E+04    4
PYRLNE    1/29/99  THERMC  4.H   5N   1    0    300.000  5000.000 1612.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 1.34940533E+01 1.30782225E-02-5.31092725E-06 9.16774974E-10-5.70507480E-14    2
 1.25447012E+04-5.29019191E+01 5.18331222E-01 3.05263735E-02-6.96325842E-06    3
-4.74435769E-09 1.85423711E-12 1.85043254E+04 2.16317664E+01                   4
PYRLYL    1/29/99  THERMC  4.H   4N   1    0    300.000  5000.000 1441.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 1.42655423E+01 7.16959055E-03-2.61629833E-06 4.24123219E-10-2.53584367E-14    2
 2.87282192E+04-5.49876875E+01-3.37777631E+00 4.89860058E-02-3.90370036E-05    3
 1.41332646E-08-1.88256423E-12 3.45930525E+04 3.92182224E+01                   4
PYROP     1/29/99  THERMC  4.H   5N   1    0    300.000  5000.000 1406.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 2.20116388E+01 2.78736506E-03-1.13805728E-06 1.97996882E-10-1.24211667E-14    2
 4.01825790E+04-9.50138981E+01-1.77243194E+01 1.29768946E-01-1.54581953E-04    3
 8.22911009E-08-1.62970458E-11 5.03953146E+04 1.05995170E+02                   4
HNCPROP   1/29/99  THERMC  4.H   5N   1    0    300.000  5000.000 1423.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 1.57166050E+01 8.54887604E-03-3.10680164E-06 5.02269358E-10-2.99741839E-14    2
 2.73052217E+04-5.90784124E+01 7.52279780E-01 3.84264182E-02-2.21149260E-05    3
 3.78397494E-09 3.31583656E-13 3.28206971E+04 2.27770410E+01                   4
A-C3H4CN  1/29/99  THERMC  4.H   4N   1    0    300.000  5000.000 1340.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 1.42039120E+01 9.92550281E-03-4.36878399E-06 7.99265452E-10-5.19044906E-14    2
 2.72109716E+04-5.18657327E+01-7.06083475E+00 6.62435950E-02-6.33711883E-05    3
 2.93828617E-08-5.33457552E-12 3.39903133E+04 6.00886287E+01                   4
C-C3H4CN  1/29/99  THERMC  4.H   4N   1    0    300.000  5000.000 1375.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 1.49368791E+01 6.47668905E-03-2.34750744E-06 3.78853855E-10-2.25817375E-14    2
 3.97271995E+04-5.00165292E+01 2.87163948E+00 3.38692899E-02-2.51401129E-05    3
 8.54475962E-09-1.06764268E-12 4.39030490E+04 1.49085502E+01                   4
C3H4CN    1/29/99  THERMC  4.H   4N   1    0    300.000  5000.000 1396.000    61 ! Martoprawiro M., Backsay G.B. & Mackie J.C., JPCA (1999) 103, 3923-3934
 1.56099688E+01 5.90248907E-03-2.14919493E-06 3.47899402E-10-2.07802288E-14    2
 3.61529551E+04-5.79376609E+01 1.63184648E+00 3.98358201E-02-3.29800298E-05    3
 1.27631797E-08-1.88643021E-12 4.07507474E+04 1.64665197E+01                   4
A-C3H5CN  1/16/17  THERMC  4.H   5N   1    2    300.000  5000.000 1430.000    61 ! Doughty, A., & Mackie, J. C., JPCA (1992) 96(1), 272-281.
 1.09928614E+01 1.45505248E-02-4.50210949E-06 6.50638889E-10-3.58287304E-14    2
 1.43674178E+04-3.11936847E+01 1.20559815E+00 4.33394942E-02-3.68365078E-05    3
 1.69025079E-08-3.09307073E-12 1.71119297E+04 1.91618447E+01                   4
T-C3H5CN  1/16/17  THERMC  4.H   5N   1    2    300.000  5000.000 1396.000    61 ! Doughty, A., & Mackie, J. C., JPCA (1992) 96(1), 272-281.
 1.09017230E+01 1.43290238E-02-5.16465461E-06 9.09557179E-10-5.91701412E-14    2
 1.16777269E+04-3.30706603E+01 1.12815965E-02 4.11350983E-02-3.09863686E-05    3
 1.24489967E-08-2.06101384E-12 1.53434572E+04 2.49667826E+01                   4
C-C3H5CN  1/16/17  THERMC  4.H   5N   1    2    300.000  5000.000 1396.000    61 ! Doughty, A., & Mackie, J. C., JPCA (1992) 96(1), 272-281.
 1.07406806E+01 1.44270533E-02-5.17031206E-06 9.06160193E-10-5.87761178E-14    2
 1.09006733E+04-3.22136921E+01-2.43844711E-01 4.14247293E-02-3.11365893E-05    3
 1.24941464E-08-2.06685041E-12 1.46026566E+04 2.63403254E+01                   4
CHCHCN CH=CHCN    A12/04C  3.H  2.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database (C3H2CN)
 6.99670220E+00 7.50618110E-03-2.68300369E-06 4.31684490E-10-2.57821318E-14    2
 5.04796219E+04-1.01552187E+01 2.15324611E+00 2.06638717E-02-1.33975241E-05    3
 7.77214839E-10 2.02897347E-12 5.18184058E+04 1.48728946E+01 5.32629680E+04    4
CH2CHCN CH2=CHCN  A12/04C  3.H  3.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database (C3H2CN)
 6.52096861E+00 1.05028771E-02-3.73734374E-06 5.99498117E-10-3.57283503E-14    2
 1.92525453E+04-9.59580896E+00 3.04396646E+00 1.05333467E-02 1.96574996E-05    3
-3.42001077E-08 1.48155667E-11 2.06456740E+04 1.05816246E+01 2.21344883E+04    4
C4H4N2 SUCCINONITRT12/03C  4.H  4.N  2.   0.G   200.000  6000.000 1000.        1
 1.14626097E+01 1.43425847E-02-5.26374167E-06 8.61140761E-10-5.20073439E-14    2
 2.02962879E+04-3.23404065E+01 2.92554100E+00 2.74517845E-02 9.39908894E-06    3
-3.65605156E-08 1.81346873E-11 2.31092217E+04 1.41181715E+01 2.52209691E+04    4
C4H3N2    1/29/99  THERMC  4.H  3.N  2.   0.G   300.000  5000.000 1537.000    61  ! K Sendt E Ikeda GB Bacskay JC Mackie JPCA 103 (1999) 1054-1072
 1.78444927E+01 5.53110368E-03-2.34526416E-06 4.17551812E-10-2.65848486E-14    2
 3.76984604E+04-6.79878141E+01 9.52114548E+00 4.46968930E-03 2.25289931E-05    3
-2.13113568E-08 5.36499501E-12 4.27060163E+04-1.58875908E+01                   4
C4H2N2    1/29/99  THERMC  4.H  2.N  2.   0.G   300.000  5000.000 1679.000    61  ! K Sendt E Ikeda GB Bacskay JC Mackie JPCA 103 (1999) 1054-1072
 1.46414829E+01 6.34973068E-03-2.73148192E-06 4.91630086E-10-3.15448650E-14    2
 3.45707689E+04-5.24954212E+01 3.10223328E+00 3.06140478E-02-2.00862591E-05    3
 5.27139118E-09-3.96461834E-13 3.86027891E+04 1.01004955E+01                   4
C2H5CN PropionitrA  1/05C  3.H  5.N  1.   0.G   200.000  6000.000 1000.        1  ! C3H5N in Burcat database
 7.04418234E+00 1.53008159E-02-5.44095595E-06 8.72156064E-10-5.19455789E-14    2
 3.05885503E+03-1.15133490E+01 3.62429314E+00 1.26256761E-02 2.47719570E-05    3
-3.99054512E-08 1.66077777E-11 4.60780029E+03 9.10669692E+00 6.39739347E+03    4
CH2CH2CN  1/29/99  THERMC  3.H  4.N  1.   0.G   300.000  5000.000 1254.000    61  ! K Sendt E Ikeda GB Bacskay JC Mackie JPCA 103 (1999) 1054-1072
 1.08023780E+01 1.04405370E-02-4.59647366E-06 8.41034552E-10-5.46218232E-14    2
 2.34914821E+04-3.44545688E+01-2.06724114E+00 3.61477061E-02-2.42081177E-05    3
 8.12552666E-09-1.22443630E-12 2.85306905E+04 3.64765218E+01                   4
CH3CHCN   1/29/99  THERMC  3.H  4.N  1.   0.G   300.000  5000.000 1681.000    61  ! K Sendt E Ikeda GB Bacskay JC Mackie JPCA 103 (1999) 1054-1072
 7.99632382E+00 1.34530512E-02-5.75498001E-06 1.03132613E-09-6.59477260E-14    2
 2.29924034E+04-1.70967993E+01 6.51512710E+00 4.37286730E-04 2.39394634E-05    3
-1.87713240E-08 4.13145742E-12 2.51173833E+04-3.19504522E+00                   4
RCTN-1   10/13/17  THERMC  4.H  6.N  1.   0.G   300.000  5000.000 1668.000    61
 1.22572997E+01 1.50342019E-02-5.63013229E-06 9.31426214E-10-5.65460201E-14    2
 2.09882388E+04-3.52340117E+01 1.61914029E+00 3.46673557E-02-1.60439742E-05    3
 1.65803319E-09 3.94529016E-13 2.49591723E+04 2.34363442E+01                   4
RCTN-2   10/13/17  THERMC  4.H  6.N  1.   0.G   300.000  5000.000 1394.000    61
 1.57305543E+01 1.05609149E-02-3.68830695E-06 5.81567945E-10-3.41348142E-14    2
 2.56241356E+04-7.38317310E+01-1.44504286E+00 4.99903036E-02-3.67034405E-05    3
 1.23812062E-08-1.51619189E-12 3.14888137E+04 1.83765220E+01                   4
ROHCTN-2 10/13/17  THERMC  4.H  6.N  1.O  1.G   300.000  5000.000 1552.000    61
 1.89520103E+01 1.10310157E-02-3.99442651E-06 6.44232539E-10-3.83826878E-14    2
 4.07565042E+03-7.87112555E+01 1.39609252E+00 4.68050754E-02-2.83676286E-05    3
 6.28313612E-09-9.63872394E-14 1.05348265E+04 1.71673874E+01                   4
RCTN-4   10/13/17  THERMC  4.H  6.N  1.   0.G   300.000  5000.000 2039.000    61
 1.35818392E+01 1.37966703E-02-5.17336426E-06 8.56608335E-10-5.20359781E-14    2
 1.51378351E+04-4.46954461E+01 1.50058258E+00 3.94849928E-02-2.39070512E-05    3
 6.22397251E-09-5.09736651E-13 1.93405098E+04 2.07418063E+01                   4
RACN-2   10/13/17  THERMC  3.H  4.N  1.   0.G   300.000  5000.000 2009.000    61
 8.53593068E+00 1.25826076E-02-5.32091919E-06 9.45696397E-10-6.01038282E-14    2
 2.67965972E+04-1.76340230E+01 6.16788913E+00 6.51532085E-03 1.28419462E-05    3
-1.18769620E-08 2.71600712E-12 2.87565365E+04-7.36582208E-01                   4
RACN-3   10/13/17  THERMC  3.H  4.N  1.   0.G   300.000  5000.000 1673.000    61
 1.91916189E+01 9.42148865E-05-4.17164564E-08 7.66087663E-12-4.99099472E-16    2
 2.56934216E+04-7.83513935E+01-1.39375456E+01 9.11267828E-02-9.36690178E-05    3
 4.27590291E-08-7.31476587E-12 3.53056414E+04 9.38719392E+01                   4
ROHACN-2 10/13/17  THERMC  3.H  4.N  1.O  1.G   300.000  5000.000 1385.000    61
 1.04261603E+01 1.44720939E-02-6.28846470E-06 1.13964934E-09-7.34834549E-14    2
 8.33074599E+03-2.60517251E+01-5.22435850E+00 6.04821849E-02-6.12785189E-05    3
 3.11780721E-08-6.15937204E-12 1.31467500E+04 5.51702242E+01                   4
ROHACN-3 10/13/17  THERMC  3.H  4.N  1.O  1.G   300.000  5000.000 1414.000    61
 1.65126224E+01 5.10968792E-03-1.86986468E-06 3.03683485E-10-1.81806834E-14    2
 8.74417336E+03-6.75145599E+01-1.24744838E-01 4.93113982E-02-4.65483707E-05    3
 2.06105205E-08-3.50635910E-12 1.38341393E+04 1.96889305E+01                   4
C4H4NO2  10/17/17  THERMC  4.H  4.N  1.O  2.G   300.000  5000.000 1396.000    61
 1.97101004E+01 7.64871349E-03-2.78308271E-06 4.50304538E-10-2.68885330E-14    2
-1.34702487E+03-7.30406448E+01 8.90040219E-01 5.48813020E-02-4.77276033E-05    3
 1.96705384E-08-3.13854266E-12 4.71031101E+03 2.66244859E+01                   4
CH2NH (H2C=NH)    T 8/11C  1.H  3.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database (CH3N)
 3.44258358E+00 8.37600036E-03-2.97819078E-06 4.77352867E-10-2.84295062E-14    2
 8.97134621E+03 3.95595397E+00 4.79302577E+00-1.26841692E-02 5.69766521E-05    3
-6.34985251E-08 2.37023330E-11 9.41385818E+03 1.10277996E+00 1.06682174E+04    4
CH2N  H2C=N*      T 1/11C  1.H  2.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat database
 3.80315578E+00 5.47197362E-03-1.95314875E-06 3.13362403E-10-1.86249384E-14    2
 2.71302747E+04 3.31759436E+00 3.97799555E+00-3.43275801E-03 2.59134260E-05    3
-3.04692171E-08 1.16272717E-11 2.74854081E+04 4.43067396E+00 2.86930920E+04    4
NCCH(3)  11/13/17  THERMC  2.H  1.N  1.   2.G   300.000  5000.000 1426.000    61
 7.05553318E+00 3.10686608E-03-2.51794650E-06 8.62579465E-10-7.93566639E-14    2
 4.30297310E+03-1.45455851E+01 3.37242258E+00 9.03135655E-03-6.11959285E-06    3
 1.99202763E-09-2.52636007E-13 6.04948556E+03 6.50451437E+00                   4
C2N   N(CC) cy    T 8/12C  2.N  1.   0.   0.G   200.000  6000.000 1000.        1
 5.31957216E+00 1.68318589E-03-6.50522050E-07 1.10121243E-10-6.80945770E-15    2
 8.53725842E+04-2.56453754E+00 3.24444516E+00 4.85727791E-03 2.60431956E-06    3
-8.16719307E-09 3.91669823E-12 8.60603450E+04 8.74664697E+00 8.72522855E+04    4
C4N2              g 6/01C  4.N  2.   0.   0.G   200.000  6000.000 1000.        1
 1.04153519E+01 5.71823954E-03-2.12579288E-06 3.50943265E-10-2.13327917E-14    2
 6.00000379E+04-2.67166250E+01 2.17476309E+00 4.76126863E-02-8.98016589E-05    3
 8.41509508E-08-2.97993323E-11 6.15242900E+04 1.16619961E+01 6.36477676E+04    4
IC4H4N2   1/14/17  THERMC  4.H  4.N  2    2.G   300.000  5000.000 1427.000    61
 1.12759705E+01 1.45352100E-02-4.54580418E-06 6.62501907E-10-3.67218596E-14    2
 2.78469747E+04-3.21423318E+01 1.56443489E+00 4.15020983E-02-3.32732837E-05    3
 1.44588523E-08-2.53553220E-12 3.07295482E+04 1.83903810E+01                   4
CH2NO                   C   1H   2N   1O   1G   200.00   6000.00 1000.00       1 !Chen, X., Fuller, M. E., & Goldsmith, C. F. React Chem Eng. (2019)
 3.87818580E+00-6.65308860E-03 5.39476100E-05-6.81768130E-08 2.71817460E-11    2
 2.57168570E+04 7.46187740E+00 5.40281520E+00 6.90570010E-03-2.51629770E-06    3
 4.10140660E-10-2.47183000E-14 2.45286900E+04-4.45742620E+00                   4
!C6H4OH                  H   5C   6O   1     G   100.000  5000.000  941.33      1 !R.D.B. New Species for Phenol
! 1.53185205E+01 1.28154562E-02-3.09306429E-06 5.36729645E-10-4.30763483E-14    2 !Species via Group / RMG.mit
! 1.30270205E+04-5.47967254E+01 1.98887816E+00 2.77378264E-02 3.96071080E-05    3 !
!-7.67853659E-08 3.29960166E-11 1.73849363E+04 1.85231300E+01                   4 !
!C6H4OH            T06/03C  6.H  5.O  1.   0.G   200.000  6000.000 1000.        1  BURCAT
! 1.29030189E+01 1.90770078E-02-6.93077391E-06 1.12768340E-09-6.78871785E-14    2
! 2.36556456E+04-4.19987250E+01 1.42119736E+00 3.09988829E-02 3.06365948E-05    3
!-6.78383584E-08 3.08907323E-11 2.77038599E+04 2.18583542E+01 2.96565883E+04    4
OOC6H4OH                H   5C   6O   3     G   100.000  5000.000  963.91      1 !R.D.B. New Species for Phenol
 1.81299995E+01 1.75612994E-02-5.77773366E-06 1.04092590E-09-7.58650187E-14    2 !Species via Group / RMG.mit
-9.94476464E+03-6.52286713E+01 7.35752801E-01 5.86569390E-02-2.13539540E-05    3 !
-2.16436322E-08 1.44851177E-11-5.14730690E+03 2.55402872E+01                   4 !
!HCCOH                   H   3C   2O   1     G   100.000  5000.000  989.31      1 !R.D.B. New Species for Phenol
! 8.13569321E+00 6.57602167E-03-2.60030811E-06 4.90280292E-10-3.53764443E-14    2 !Species via RMG.mit : Source: Klippenstein
! 1.30908011E+04-1.75941492E+01 3.01766475E+00 1.74503768E-02-4.20053610E-06    3 !
!-8.46362785E-09 4.76244533E-12 1.45839741E+04 9.47087842E+00                   4 !
!OHBENZYNE               H   4C   6O   1     G   100.000  5000.000  961.91      1 !R.D.B. New Species for Phenol
! 1.57981076E+01 1.14731374E-02-3.60923434E-06 6.83108180E-10-5.30527141E-14    2 !Species via Group / RMG.mit
! 2.37538903E+04-5.96871714E+01 1.63018169E+00 3.93376946E-02 1.36010369E-06    3 !
!-3.63200859E-08 1.82860653E-11 2.79160844E+04 1.55818037E+01                   4 !
!C6H3O2                  H   3C   6O   2     G   100.000  5000.000  988.62      1 !R.D.B. New Species for Phenol
! 1.34120746E+01 1.79858046E-02-7.48346248E-06 1.41065636E-09-1.00527990E-13    2 !Species via Group / RMG.mit / Currane Pentane
! 1.13762200E+04-4.27445680E+01 1.63426611E+00 4.19756724E-02-7.97810014E-06    3 !
!-2.24677796E-08 1.20605222E-11 1.48613728E+04 1.97903178E+01                   4 !   
FC10H10                 C  10H  10          G    300.00   4000.00 2043.00      1
 .196465049E+02 .362867673E-01-.135117921E-04 .222712581E-08-.134868100E-12    2
 .466515480E+04-.883925826E+02-.975555457E+01 .989343734E-01-.593843991E-04    3
 .154882804E-07-.129445409E-11 .148791325E+05 .708155586E+02                   4
PROTC                   C 500H 450O  65N  80S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
PROTH                                       S    300.00   5000.00 1000.00      1&
    C  400   H     900    O 150  N  86      
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
PROTO                   C 250H 500O 200N  72S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
GNH3NO                  C   0H   3O   1N   2S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
PROTOH                  C  45H  70O  25N  10S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
PROTCC                  C  90H  70O   3N  15S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
NH3S                    H   3N   1          S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
HCNS                    C   1H   1N   1     S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
CHARN                   N   1               S    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
TARN                    C  13H  15O   3N   4G    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
NH3                     H   3N   1          G    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
NO                      C   0H   0O   1N   1G    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
HCN                     C   1H   1N   1     G    300.00   5000.00 1000.00      1
 .299142300E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033800E+03-.135511000E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
C6H6                    C   6H   6          G    300.00   4000.00 1000.00      1! Burcat kik
 1.10809576E+01 2.07176746E-02-7.52145991E-06 1.22320984E-09-7.36091279E-14    2
 4.30641035E+03-4.00413310E+01 5.04818632E-01 1.85020642E-02 7.38345881E-05    3
-1.18135741E-07 5.07210429E-11 8.55247913E+03 2.16412893E+01 9.96811598E+03    4   
CELL                    C   6H  10O   5     S 300.0    4000.0    1000.0        1
 2.92532475e+01 1.95021650e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.22499447e+05 0.00000000e+00 2.92532475e+01 1.95021650e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.22499447e+05 0.00000000e+00                   4
GMSW                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38359995e+01 1.58906663e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.03125432e+05 0.00000000e+00 2.38359995e+01 1.58906663e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.03125432e+05 0.00000000e+00                   4
XYHW                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38359995e+01 1.58906663e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.07190349e+05 0.00000000e+00 2.38359995e+01 1.58906663e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.07190349e+05 0.00000000e+00                   4
XYGR                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38359995e+01 1.58906663e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.09860883e+05 0.00000000e+00 2.38359995e+01 1.58906663e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.09860883e+05 0.00000000e+00                   4
LIGC                    C  15H  14O   4     S 300.0    4000.0    1000.0        1
 4.65972456e+01 3.10648304e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.01283047e+05 0.00000000e+00 4.65972456e+01 3.10648304e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.01283047e+05 0.00000000e+00                   4
LIGH                    C  22H  28O   9     S 300.0    4000.0    1000.0        1
 7.87449483e+01 5.24966322e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.23767540e+05 0.00000000e+00 7.87449483e+01 5.24966322e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.23767540e+05 0.00000000e+00                   4
LIGO                    C  20H  22O  10     S 300.0    4000.0    1000.0        1
 7.62062786e+01 5.08041857e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.51431603e+05 0.00000000e+00 7.62062786e+01 5.08041857e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.51431603e+05 0.00000000e+00                   4
TGL                     C  57H 100O   7     S 300.0    4000.0    1000.0        1
 1.61911234e+02 1.07940823e-01 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.44639069e+05 0.00000000e+00 1.61911234e+02 1.07940823e-01 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.44639069e+05 0.00000000e+00                   4
TANN                    C  15H  12O   7     S 300.0    4000.0    1000.0        1
 5.48930719e+01 3.65953813e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.60348491e+05 0.00000000e+00 5.48930719e+01 3.65953813e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.60348491e+05 0.00000000e+00                   4
TANNH                   C   8H   6O   5     S 300.0    4000.0    1000.0        1
 5.48900197e+01 3.65933465e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.59515809e+05 0.00000000e+00 5.48900197e+01 3.65933465e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.59515809e+05 0.00000000e+00                   4 !!!MUST SET THE PARAMETERS CORRECTLY
!MOIST                   C   0H   2O   1     S 300.0    4000.0    1000.0        1   !From DH vaporization  engineering tool box
! 9.04470000E+00 1.60000000E-03-6.00000000E-06 6.00000000E-09-2.00000000E-12    2
!-3.70865499E+04-2.88280137E+02 9.04470000E+00 1.60000000E-03-6.00000000E-06    3
! 6.00000000E-09-2.00000000E-12-3.70865499E+04-2.88280137E+02                   4
MOIST                   C   0H   2O   1     S 300.0    4000.0    1000.0        1   !LOW T FROM BURCAT. HIGH T FROM DHR
 3.25005985e+00 2.16670657e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-3.49947368e+04 0.00000000e+00 7.25575005E+01-6.62445402E-01 2.56198746E-03    3
-4.36591923E-06 2.78178981E-09-4.18865499E+04-2.88280137E+02                   4
ASH                     C   0H   0K   1     S 300.0    4000.0    1000.0        1
 7.05472697e+00 4.70315131e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-6.09058102e+03 0.00000000e+00 7.05472697e+00 4.70315131e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-6.09058102e+03 0.00000000e+00                   4
CELLA                   C   6H  10O   5     S 300.0    4000.0    1000.0        1
 2.92532475e+01 1.95021650e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25202436e+05 0.00000000e+00 2.92532475e+01 1.95021650e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25202436e+05 0.00000000e+00                   4
HCE1                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38359995e+01 1.58906663e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.92805242e+04 0.00000000e+00 2.38359995e+01 1.58906663e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.92805242e+04 0.00000000e+00                   4
HCE2                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38359995e+01 1.58906663e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.10893282e+05 0.00000000e+00 2.38359995e+01 1.58906663e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.10893282e+05 0.00000000e+00                   4
LIGCC                   C  15H  14O   4     S 300.0    4000.0    1000.0        1
 4.65972456e+01 3.10648304e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-7.01136192e+04 0.00000000e+00 4.65972456e+01 3.10648304e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-7.01136192e+04 0.00000000e+00                   4
LIGOH                   C  19H  22O   8     S 300.0    4000.0    1000.0        1
 6.82662377e+01 4.55108251e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.86155940e+05 0.00000000e+00 6.82662377e+01 4.55108251e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.86155940e+05 0.00000000e+00                   4
LIG                     C  11H  12O   4     S 300.0    4000.0    1000.0        1
 3.75654919e+01 2.50436613e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.43494885e+04 0.00000000e+00 3.75654919e+01 2.50436613e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.43494885e+04 0.00000000e+00                   4
ITANN                   C   8H   4O   4     S 300.0    4000.0    1000.0        1
 5.48930719e+01 3.65953813e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.60348491e+05 0.00000000e+00 5.48930719e+01 3.65953813e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.60348491e+05 0.00000000e+00                   4
CHAR                    C   1               S 300.0    4000.0    1000.0        1
-1.00801964e-01 4.99856387e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-4.20593720e+02 0.00000000e+00-1.00801964e-01 4.99856387e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-4.20593720e+02 0.00000000e+00                   4
CHARO                   C   1H   0O   1     S 300.0    4000.0    1000.0        1
-2.35073100e-01 1.16567958e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.47486517e+03 0.00000000e+00-2.35073100e-01 1.16567958e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.47486517e+03 0.00000000e+00                   4
COH2S                   C   1H   2O   1     S 300.0    4000.0    1000.0        1
 5.41724802e+00 3.61149868e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-4.29716079e+04 0.00000000e+00 5.41724802e+00 3.61149868e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-4.29716079e+04 0.00000000e+00                   4
CO2S                    C   1H   0O   2     S 300.0    4000.0    1000.0        1
 7.94004089e+00 5.29336060e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-3.99924651e+04 0.00000000e+00 7.94004089e+00 5.29336060e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-3.99924651e+04 0.00000000e+00                   4
COS                     C   1H   0O   1     S 300.0    4000.0    1000.0        1
 5.05352418e+00 3.36901612e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.01008627e+04 0.00000000e+00 5.05352418e+00 3.36901612e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.01008627e+04 0.00000000e+00                   4
COSTIFFS                C   1H   0O   1     S 300.0    4000.0    1000.0        1
 5.05352418e+00 3.36901612e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.46120426e+03 0.00000000e+00 5.05352418e+00 3.36901612e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.46120426e+03 0.00000000e+00                   4
CH3OHS                  C   1H   4O   1     S 300.0    4000.0    1000.0        1
 5.78097185e+00 3.85398124e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.62398341e+04 0.00000000e+00 5.78097185e+00 3.85398124e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.62398341e+04 0.00000000e+00                   4
CH4S                    C   1H   4O   0     S 300.0    4000.0    1000.0        1
 2.89445514e+00 1.92963676e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.10504531e+03 0.00000000e+00 2.89445514e+00 1.92963676e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.10504531e+03 0.00000000e+00                   4
C2H4S                   C   2H   4O   0     S 300.0    4000.0    1000.0        1
 5.06146259e+00 3.37430840e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
 5.04456594e+03 0.00000000e+00 5.06146259e+00 3.37430840e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00 5.04456594e+03 0.00000000e+00                   4
C6H5OHS                 C   6H   6O   1     S 300.0    4000.0    1000.0        1
 1.69797330e+01 1.13198220e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.86147802e+04 0.00000000e+00 1.69797330e+01 1.13198220e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.86147802e+04 0.00000000e+00                   4
CH2OS                   C   1H   2O   1     S 300.0    4000.0    1000.0        1
 5.41724802e+00 3.61149868e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.46988983e+04 0.00000000e+00 5.41724802e+00 3.61149868e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.46988983e+04 0.00000000e+00                   4
H2S                     C   0H   2O   0     S 300.0    4000.0    1000.0        1
 3.63723839e-01 2.42482560e-04 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
 7.83252454e+02 0.00000000e+00 3.63723839e-01 2.42482560e-04 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00 7.83252454e+02 0.00000000e+00                   4
C2H6S                   C   2H   6O   0     S 300.0    4000.0    1000.0        1
 5.42518643e+00 3.61679096e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.10383524e+04 0.00000000e+00 5.42518643e+00 3.61679096e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.10383524e+04 0.00000000e+00                   4
VANILLIN                C   8H   8O   3     G    300.00   3500.00 1260.00      1
 1.36544650e+01 4.84143232e-02-2.42641798e-05 5.50487829e-09-4.76001947e-13    2
-5.18855416e+04-3.54575728e+01-4.86637458e+00 1.07210639e-01-9.42597942e-05    3
 4.25395949e-08-7.82416000e-12-4.72182900e+04 5.81751551e+01                   4
CRESOL                  C   7H   8O   1     G    300.00   4000.00 1000.00      1
 .109411883E+02 .359221340E-01-.155859930E-04 .305336930E-08-.221926260E-12    2
-.211837368E+05-.322120090E+02-.410479790E+01 .823735850E-01-.680002460E-04    3
 .287114670E-07-.487123580E-11-.173767210E+05 .440872850E+02                   4
LVGS                    C   6H  10O   5     S 300.0    4000.0    1000.0        1
 2.92532475e+01 1.95021650e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25616758e+05 0.00000000e+00 2.92532475e+01 1.95021650e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25616758e+05 0.00000000e+00                   4
END
