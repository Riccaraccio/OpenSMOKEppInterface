   THERMO 
   300.0   1000.0   3000.0
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2
-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3
 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00 0.00000000E+00    4
BIOMASS                 C   6H  10O   5     S 300.0    4000.0    1000.0        1!From CELL
 2.92516210e+01 1.95010807e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25919988e+05 0.00000000e+00 2.92516210e+01 1.95010807e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25919988e+05 0.00000000e+00                   4
H2O               ATcT3EH   2O   1    0    0G    200.00   6000.00 1000.00      1
 2.73117512E+00 2.95136995E-03-8.35359785E-07 1.26088593E-10-8.40531676E-15    2
-2.99169082E+04 6.55183000E+00 4.20147551E+00-2.05583546E-03 6.56547207E-06    3
-5.52906960E-09 1.78282605E-12-3.02950066E+04-8.60610906E-01-2.90858262E+04    4
CHAR                    C   1               S 300.0    4000.0    1000.0        1
-1.00796361E-01	4.99828606E-03 0.00000000E+00 0.00000000E+00 0.00000000E+00    2           
-1.94683964E+02 0.00000000E+00-1.00796361E-01 4.99828606E-03 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.94683964E+02 0.00000000E+00                   4
TAR                     C   6H  10O   5     S 300.0    4000.0    1000.0        1!From CELL
 .279850422E+02 .264166682E-01-.913640739E-05 .142923991E-08-.833656585E-13    2
-.114313686E+06-.117754445E+03-.781241700E+01 .125424511E+00-.116271866E-03    3
 .544734561E-07-.100746170E-10-.103428291E+06 .690300863E+02                   4
CO                ATcT3EC   1O   1    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] CO <g> ATcT ver. 1.122, DHf298 = -110.523 � 0.026 kJ/mol - fit MAR17
 3.03397274E+00 1.37328118E-03-4.96445087E-07 8.10281447E-11-4.85331749E-15    2
-1.42586044E+04 6.10076092E+00 3.59508377E+00-7.21196937E-04 1.28238234E-06    3
 6.52429293E-10-8.21714806E-13-1.43448968E+04 3.44355598E+00-1.32928623E+04    4
CO2               ATcT3EC   1O   2    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] CO2 <g> ATcT ver. 1.122, DHf298 = -393.475 � 0.015 kJ/mol - fit MAR17
 4.63537470E+00 2.74559459E-03-9.98282389E-07 1.61013606E-10-9.22018642E-15    2
-4.90203677E+04-1.92887630E+00 2.20664321E+00 1.00970086E-02-9.96338809E-06    3
 5.47155623E-09-1.27733965E-12-4.83529864E+04 1.05261943E+01-4.73241678E+04    4
O2                ATcT3EO   2    0    0    0G    200.00   6000.00 1000.00      1	! [Ghobad] O2 <g> ATcT ver. 1.122, DHf298 = 0.000 � 0.000 kJ/mol - fit MAR17
 3.65980488E+00 6.59877372E-04-1.44158172E-07 2.14656037E-11-1.36503784E-15    2
-1.21603048E+03 3.42074148E+00 3.78498258E+00-3.02002233E-03 9.92029171E-06    3
-9.77840434E-09 3.28877702E-12-1.06413589E+03 3.64780709E+00 0.00000000E+00    4
CH4               G 8/99C  1 H  4    0    0 G   200.000  6000.00  1000.00      1
 1.65326226E+00 1.00263099E-02-3.31661238E-06 5.36483138E-10-3.14696758E-14    2
-1.00095936E+04 9.90506283E+00 5.14911468E+00-1.36622009E-02 4.91453921E-05    3
-4.84246767E-08 1.66603441E-11-1.02465983E+04-4.63848842E+00-8.97226656E+03    4
H2                ATcT3EH   2    0    0    0G    200.00   6000.00 1000.00      1
 2.90207649E+00 8.68992581E-04-1.65864430E-07 1.90851899E-11-9.31121789E-16    2
-7.97948726E+02-8.45591320E-01 2.37694204E+00 7.73916922E-03-1.88735073E-05    3
 1.95517114E-08-7.17095663E-12-9.21173081E+02 5.47184736E-01 0.00000000E+00    4
MOIST                   C   0H   2O   1     S 300.0    4000.0    1000.0        1
 3.25005985e+00 2.16670657e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-3.49947368e+04 0.00000000e+00 7.25575005E+01-6.62445402E-01 2.56198746E-03    3
-4.36591923E-06 2.78178981E-09-4.18865499E+04-2.88280137E+02                   4
